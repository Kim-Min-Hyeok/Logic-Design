<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-59.2333,11.6667,126.633,-81.8</PageViewport>
<gate>
<ID>2</ID>
<type>AE_FULLADDER_4BIT</type>
<position>81,-22.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>10 </input>
<input>
<ID>IN_3</ID>9 </input>
<input>
<ID>IN_B_0</ID>16 </input>
<input>
<ID>IN_B_1</ID>15 </input>
<input>
<ID>IN_B_2</ID>14 </input>
<input>
<ID>IN_B_3</ID>13 </input>
<output>
<ID>OUT_0</ID>26 </output>
<output>
<ID>OUT_1</ID>19 </output>
<output>
<ID>OUT_2</ID>22 </output>
<output>
<ID>OUT_3</ID>20 </output>
<input>
<ID>carry_in</ID>17 </input>
<output>
<ID>carry_out</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>4</ID>
<type>AE_FULLADDER_4BIT</type>
<position>7.5,-22.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>2 </input>
<input>
<ID>IN_3</ID>1 </input>
<input>
<ID>IN_B_0</ID>8 </input>
<input>
<ID>IN_B_1</ID>7 </input>
<input>
<ID>IN_B_2</ID>6 </input>
<input>
<ID>IN_B_3</ID>5 </input>
<output>
<ID>OUT_0</ID>40 </output>
<output>
<ID>OUT_1</ID>38 </output>
<output>
<ID>OUT_2</ID>39 </output>
<output>
<ID>OUT_3</ID>34 </output>
<input>
<ID>carry_in</ID>25 </input>
<output>
<ID>carry_out</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>-0.5,-16</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>-0.5,-12.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>-0.5,-9</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>-0.5,-5.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>7,-16</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>7,-12.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>7,-9</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>7,-5.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>73.5,-16</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>73.5,-12.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>73.5,-9</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>73.5,-5.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>80.5,-5.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>80.5,-9</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>80.5,-12.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>80.5,-16</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>87.5,-16</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>AE_FULLADDER_4BIT</type>
<position>77.5,-38</position>
<input>
<ID>IN_1</ID>25 </input>
<input>
<ID>IN_2</ID>25 </input>
<input>
<ID>IN_B_0</ID>26 </input>
<input>
<ID>IN_B_1</ID>19 </input>
<input>
<ID>IN_B_2</ID>22 </input>
<input>
<ID>IN_B_3</ID>20 </input>
<output>
<ID>OUT_0</ID>27 </output>
<output>
<ID>OUT_1</ID>30 </output>
<output>
<ID>OUT_2</ID>31 </output>
<output>
<ID>OUT_3</ID>33 </output>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>50</ID>
<type>AE_FULLADDER_4BIT</type>
<position>4,-38</position>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>41 </input>
<input>
<ID>IN_B_0</ID>40 </input>
<input>
<ID>IN_B_1</ID>38 </input>
<input>
<ID>IN_B_2</ID>39 </input>
<input>
<ID>IN_B_3</ID>34 </input>
<output>
<ID>OUT_0</ID>46 </output>
<output>
<ID>OUT_1</ID>44 </output>
<output>
<ID>OUT_2</ID>43 </output>
<output>
<ID>OUT_3</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>54</ID>
<type>AE_OR3</type>
<position>123.5,-17</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>23 </input>
<input>
<ID>IN_2</ID>24 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_AND2</type>
<position>110.5,-17</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_AND2</type>
<position>110.5,-22.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>GA_LED</type>
<position>82,-44.5</position>
<input>
<ID>N_in3</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>79,-44.5</position>
<input>
<ID>N_in3</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>GA_LED</type>
<position>76,-44.5</position>
<input>
<ID>N_in3</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>GA_LED</type>
<position>73,-44.5</position>
<input>
<ID>N_in3</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AE_OR3</type>
<position>54.5,-17</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>35 </input>
<input>
<ID>IN_2</ID>36 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND2</type>
<position>40,-17</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_AND2</type>
<position>40,-22.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>GA_LED</type>
<position>5.5,-44.5</position>
<input>
<ID>N_in3</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>GA_LED</type>
<position>8.5,-44.5</position>
<input>
<ID>N_in3</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>GA_LED</type>
<position>2.5,-44.5</position>
<input>
<ID>N_in3</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>GA_LED</type>
<position>-0.5,-44.5</position>
<input>
<ID>N_in3</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>-9,-44.5</position>
<input>
<ID>N_in3</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>82.5,-0.5</position>
<gparam>LABEL_TEXT B1's</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>75,-0.5</position>
<gparam>LABEL_TEXT A1's</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>9,-1.5</position>
<gparam>LABEL_TEXT B2's</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>1,-1.5</position>
<gparam>LABEL_TEXT A2's</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>-9.5,-47</position>
<gparam>LABEL_TEXT Cout</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_LABEL</type>
<position>3.5,-47</position>
<gparam>LABEL_TEXT sum2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>77.5,-47</position>
<gparam>LABEL_TEXT sum1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-18.5,2.5,-16</points>
<connection>
<GID>4</GID>
<name>IN_3</name></connection>
<intersection>-16 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>1.5,-16,2.5,-16</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-18.5,3.5,-12.5</points>
<connection>
<GID>4</GID>
<name>IN_2</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1.5,-12.5,3.5,-12.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-18.5,4.5,-9</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1.5,-9,4.5,-9</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-18.5,5.5,-5.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1.5,-5.5,5.5,-5.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9.5,-18.5,9.5,-16</points>
<connection>
<GID>4</GID>
<name>IN_B_3</name></connection>
<intersection>-16 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>9,-16,9.5,-16</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-18.5,10.5,-12.5</points>
<connection>
<GID>4</GID>
<name>IN_B_2</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-12.5,10.5,-12.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11.5,-18.5,11.5,-9</points>
<connection>
<GID>4</GID>
<name>IN_B_1</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-9,11.5,-9</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-18.5,12.5,-5.5</points>
<connection>
<GID>4</GID>
<name>IN_B_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-5.5,12.5,-5.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-18.5,76,-16</points>
<connection>
<GID>2</GID>
<name>IN_3</name></connection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>75.5,-16,76,-16</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-18.5,77,-12.5</points>
<connection>
<GID>2</GID>
<name>IN_2</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-12.5,77,-12.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-18.5,78,-9</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-9,78,-9</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-18.5,79,-5.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-5.5,79,-5.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-18.5,83,-16</points>
<connection>
<GID>2</GID>
<name>IN_B_3</name></connection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-16,83,-16</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-18.5,84,-12.5</points>
<connection>
<GID>2</GID>
<name>IN_B_2</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-12.5,84,-12.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-18.5,85,-9</points>
<connection>
<GID>2</GID>
<name>IN_B_1</name></connection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-9,85,-9</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-18.5,86,-5.5</points>
<connection>
<GID>2</GID>
<name>IN_B_0</name></connection>
<intersection>-5.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-5.5,86,-5.5</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-21.5,89.5,-16</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89,-21.5,89.5,-21.5</points>
<connection>
<GID>2</GID>
<name>carry_in</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81.5,-27,96.5,-27</points>
<intersection>81.5 4</intersection>
<intersection>81.5 4</intersection>
<intersection>96.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>96.5,-27,96.5,-16</points>
<intersection>-27 1</intersection>
<intersection>-16 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>96.5,-16,107.5,-16</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>96.5 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>81.5,-34,81.5,-26.5</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<connection>
<GID>48</GID>
<name>IN_B_1</name></connection>
<intersection>-27 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-34,79.5,-26.5</points>
<connection>
<GID>48</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79.5,-28,98,-28</points>
<intersection>79.5 0</intersection>
<intersection>98 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>98,-28,98,-18</points>
<intersection>-28 1</intersection>
<intersection>-18 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>98,-18,107.5,-18</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>98 2</intersection>
<intersection>103.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>103.5,-23.5,103.5,-18</points>
<intersection>-23.5 5</intersection>
<intersection>-18 3</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>103.5,-23.5,107.5,-23.5</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>103.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-2.5,120,-2.5</points>
<intersection>70 3</intersection>
<intersection>120 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70,-21.5,70,-2.5</points>
<intersection>-21.5 4</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>70,-21.5,73,-21.5</points>
<connection>
<GID>2</GID>
<name>carry_out</name></connection>
<intersection>70 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>120,-15,120,-2.5</points>
<intersection>-15 6</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>120,-15,120.5,-15</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>120 5</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-34,80.5,-26.5</points>
<connection>
<GID>48</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-29,99.5,-29</points>
<intersection>80.5 0</intersection>
<intersection>99.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>99.5,-29,99.5,-21.5</points>
<intersection>-29 1</intersection>
<intersection>-21.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>99.5,-21.5,107.5,-21.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>99.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>113.5,-17,120.5,-17</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<connection>
<GID>54</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-22.5,116.5,-19</points>
<intersection>-22.5 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-19,120.5,-19</points>
<connection>
<GID>54</GID>
<name>IN_2</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-22.5,116.5,-22.5</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-32,67,3</points>
<intersection>-32 1</intersection>
<intersection>3 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-32,126.5,-32</points>
<intersection>67 0</intersection>
<intersection>73.5 8</intersection>
<intersection>74.5 4</intersection>
<intersection>126.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>126.5,-32,126.5,-17</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>74.5,-34,74.5,-32</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>15.5,3,67,3</points>
<intersection>15.5 10</intersection>
<intersection>67 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>73.5,-34,73.5,-32</points>
<connection>
<GID>48</GID>
<name>IN_2</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>15.5,-21.5,15.5,3</points>
<connection>
<GID>4</GID>
<name>carry_in</name></connection>
<intersection>3 5</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-34,82.5,-26.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<connection>
<GID>48</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-43.5,82,-42</points>
<connection>
<GID>60</GID>
<name>N_in3</name></connection>
<intersection>-42 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>79,-42,82,-42</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>82 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-43.5,79,-42.5</points>
<connection>
<GID>62</GID>
<name>N_in3</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>78,-42.5,78,-42</points>
<connection>
<GID>48</GID>
<name>OUT_1</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>78,-42.5,79,-42.5</points>
<intersection>78 1</intersection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-43.5,76,-42.5</points>
<connection>
<GID>66</GID>
<name>N_in3</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>77,-42.5,77,-42</points>
<connection>
<GID>48</GID>
<name>OUT_2</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>76,-42.5,77,-42.5</points>
<intersection>76 0</intersection>
<intersection>77 1</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-43.5,73,-42</points>
<connection>
<GID>68</GID>
<name>N_in3</name></connection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>73,-42,76,-42</points>
<connection>
<GID>48</GID>
<name>OUT_3</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>25,-18,37,-18</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>25 4</intersection>
<intersection>31.5 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>25,-28,25,-18</points>
<intersection>-28 6</intersection>
<intersection>-18 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>6,-28,25,-28</points>
<intersection>6 7</intersection>
<intersection>6 7</intersection>
<intersection>25 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>6,-34,6,-26.5</points>
<connection>
<GID>4</GID>
<name>OUT_3</name></connection>
<connection>
<GID>50</GID>
<name>IN_B_3</name></connection>
<intersection>-28 6</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>31.5,-23.5,31.5,-18</points>
<intersection>-23.5 9</intersection>
<intersection>-18 3</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>31.5,-23.5,37,-23.5</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>31.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>43,-17,51.5,-17</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<connection>
<GID>70</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-22.5,46,-19</points>
<intersection>-22.5 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46,-19,51.5,-19</points>
<connection>
<GID>69</GID>
<name>IN_2</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-22.5,46,-22.5</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4,-0.5,51.5,-0.5</points>
<intersection>-4 15</intersection>
<intersection>51.5 16</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-4,-21.5,-4,-0.5</points>
<intersection>-21.5 17</intersection>
<intersection>-0.5 1</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>51.5,-15,51.5,-0.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>-4,-21.5,-0.5,-21.5</points>
<connection>
<GID>4</GID>
<name>carry_out</name></connection>
<intersection>-4 15</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-34,8,-26.5</points>
<connection>
<GID>50</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>4</GID>
<name>OUT_1</name></connection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-27,23.5,-27</points>
<intersection>8 0</intersection>
<intersection>23.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>23.5,-27,23.5,-16</points>
<intersection>-27 1</intersection>
<intersection>-16 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>23.5,-16,37,-16</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>23.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-34,7,-26.5</points>
<connection>
<GID>50</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>4</GID>
<name>OUT_2</name></connection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7,-29,26.5,-29</points>
<intersection>7 0</intersection>
<intersection>26.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>26.5,-29,26.5,-21.5</points>
<intersection>-29 1</intersection>
<intersection>-21.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>26.5,-21.5,37,-21.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>26.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-34,9,-26.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<connection>
<GID>50</GID>
<name>IN_B_0</name></connection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-34,0,-32</points>
<connection>
<GID>50</GID>
<name>IN_2</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9,-32,57.5,-32</points>
<intersection>-9 6</intersection>
<intersection>0 0</intersection>
<intersection>1 4</intersection>
<intersection>57.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>57.5,-32,57.5,-17</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>1,-34,1,-32</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-9,-43.5,-9,-32</points>
<connection>
<GID>81</GID>
<name>N_in3</name></connection>
<intersection>-32 1</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-43.5,-0.5,-42</points>
<connection>
<GID>79</GID>
<name>N_in3</name></connection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,-42,2.5,-42</points>
<connection>
<GID>50</GID>
<name>OUT_3</name></connection>
<intersection>-0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-42.5,3.5,-42</points>
<connection>
<GID>50</GID>
<name>OUT_2</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>2.5,-43.5,2.5,-42.5</points>
<connection>
<GID>77</GID>
<name>N_in3</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>2.5,-42.5,3.5,-42.5</points>
<intersection>2.5 1</intersection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-42.5,4.5,-42</points>
<connection>
<GID>50</GID>
<name>OUT_1</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>5.5,-43.5,5.5,-42.5</points>
<connection>
<GID>73</GID>
<name>N_in3</name></connection>
<intersection>-42.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-42.5,5.5,-42.5</points>
<intersection>4.5 0</intersection>
<intersection>5.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>8.5,-43.5,8.5,-42</points>
<connection>
<GID>75</GID>
<name>N_in3</name></connection>
<intersection>-42 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>5.5,-42,8.5,-42</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>8.5 1</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 9></circuit>