<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-23.2333,11.6667,35.7,-49.8</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>37.5,-32</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2</ID>
<type>GA_LED</type>
<position>43.5,-51</position>
<input>
<ID>N_in2</ID>1 </input>
<input>
<ID>N_in3</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>GA_LED</type>
<position>65,-51</position>
<input>
<ID>N_in2</ID>2 </input>
<input>
<ID>N_in3</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>GA_LED</type>
<position>86,-51</position>
<input>
<ID>N_in2</ID>3 </input>
<input>
<ID>N_in3</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>GA_LED</type>
<position>103,-50.5</position>
<input>
<ID>N_in2</ID>13 </input>
<input>
<ID>N_in3</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AE_DFF_LOW</type>
<position>132,-40</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>31 </output>
<input>
<ID>clock</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7</ID>
<type>GA_LED</type>
<position>142,-51</position>
<input>
<ID>N_in2</ID>4 </input>
<input>
<ID>N_in3</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AE_DFF_LOW</type>
<position>114,-40</position>
<input>
<ID>IN_0</ID>35 </input>
<output>
<ID>OUT_0</ID>32 </output>
<input>
<ID>clock</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>9</ID>
<type>GA_LED</type>
<position>124.5,-51</position>
<input>
<ID>N_in2</ID>14 </input>
<input>
<ID>N_in3</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>108,-24</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_AND3</type>
<position>114.5,-24</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>15 </input>
<input>
<ID>IN_2</ID>5 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_OR2</type>
<position>111.5,-30.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_AND2</type>
<position>25,-24</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>30.5,-24</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_AND3</type>
<position>37,-24</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>2 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_OR3</type>
<position>30.5,-30.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>36 </input>
<input>
<ID>IN_2</ID>37 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_AND2</type>
<position>46.5,-24</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>52,-24</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_AND3</type>
<position>58.5,-24</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<input>
<ID>IN_2</ID>7 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_SMALL_INVERTER</type>
<position>33.5,-10</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>21</ID>
<type>AE_SMALL_INVERTER</type>
<position>38.5,-10</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_SMALL_INVERTER</type>
<position>43.5,-10</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>23</ID>
<type>AE_SMALL_INVERTER</type>
<position>48,-10</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_SMALL_INVERTER</type>
<position>52.5,-10</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_SMALL_INVERTER</type>
<position>57,-10</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_OR3</type>
<position>52,-30.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>8 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_AND2</type>
<position>68,-24</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_AND3</type>
<position>74.5,-24</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>13 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>29</ID>
<type>AE_OR2</type>
<position>71.5,-30.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND2</type>
<position>84,-24</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_AND2</type>
<position>89.5,-24</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_AND4</type>
<position>97,-24</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>16 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>33</ID>
<type>AE_OR3</type>
<position>89.5,-30.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>18 </input>
<input>
<ID>IN_2</ID>20 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>34</ID>
<type>AE_DFF_LOW</type>
<position>37.5,-40</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>27 </output>
<input>
<ID>clear</ID>26 </input>
<input>
<ID>clock</ID>24 </input>
<input>
<ID>set</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>35</ID>
<type>AE_DFF_LOW</type>
<position>57.5,-40</position>
<input>
<ID>IN_0</ID>21 </input>
<output>
<ID>OUT_0</ID>28 </output>
<input>
<ID>clear</ID>26 </input>
<input>
<ID>clock</ID>24 </input>
<input>
<ID>set</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>36</ID>
<type>AE_DFF_LOW</type>
<position>77,-40</position>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>29 </output>
<input>
<ID>clear</ID>26 </input>
<input>
<ID>clock</ID>24 </input>
<input>
<ID>set</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>37</ID>
<type>AE_DFF_LOW</type>
<position>96,-40</position>
<input>
<ID>IN_0</ID>23 </input>
<output>
<ID>OUT_0</ID>30 </output>
<input>
<ID>clear</ID>26 </input>
<input>
<ID>clock</ID>24 </input>
<input>
<ID>set</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>37.5,-47.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>BB_CLOCK</type>
<position>26,-41</position>
<output>
<ID>CLK</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-52.5,16.5,-8</points>
<intersection>-52.5 9</intersection>
<intersection>-8 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>16.5,-8,33.5,-8</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>16.5 0</intersection>
<intersection>24 12</intersection>
<intersection>29.5 14</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>16.5,-52.5,43.5,-52.5</points>
<intersection>16.5 0</intersection>
<intersection>43.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>43.5,-52.5,43.5,-52</points>
<connection>
<GID>2</GID>
<name>N_in2</name></connection>
<intersection>-52.5 9</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>24,-21,24,-8</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>-8 7</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>29.5,-21,29.5,-8</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-8 7</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-54.5,36,-8</points>
<intersection>-54.5 13</intersection>
<intersection>-20 3</intersection>
<intersection>-8 23</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>35,-20,51,-20</points>
<intersection>35 20</intersection>
<intersection>36 0</intersection>
<intersection>45.5 4</intersection>
<intersection>51 17</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>45.5,-21,45.5,-20</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>-20 3</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>36,-54.5,65,-54.5</points>
<intersection>36 0</intersection>
<intersection>65 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>65,-54.5,65,-52</points>
<connection>
<GID>3</GID>
<name>N_in2</name></connection>
<intersection>-54.5 13</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>51,-21,51,-20</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>-20 3</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>35,-21,35,-20</points>
<connection>
<GID>15</GID>
<name>IN_2</name></connection>
<intersection>-20 3</intersection></vsegment>
<hsegment>
<ID>23</ID>
<points>36,-8,38.5,-8</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-56.5,41,-8</points>
<intersection>-56.5 16</intersection>
<intersection>-20.5 18</intersection>
<intersection>-18 8</intersection>
<intersection>-8 10</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>41,-18,58.5,-18</points>
<intersection>41 0</intersection>
<intersection>58.5 12</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>41,-8,43.5,-8</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>41 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>58.5,-21,58.5,-18</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>-18 8</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>41,-56.5,86,-56.5</points>
<intersection>41 0</intersection>
<intersection>86 17</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>86,-56.5,86,-52</points>
<connection>
<GID>4</GID>
<name>N_in2</name></connection>
<intersection>-56.5 16</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>37,-20.5,67,-20.5</points>
<intersection>37 23</intersection>
<intersection>41 0</intersection>
<intersection>67 21</intersection></hsegment>
<vsegment>
<ID>21</ID>
<points>67,-21,67,-20.5</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>-20.5 18</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>37,-21,37,-20.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>-20.5 18</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>54.5,-62.5,54.5,-8</points>
<intersection>-62.5 17</intersection>
<intersection>-21 19</intersection>
<intersection>-19.5 2</intersection>
<intersection>-8 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-19.5,100,-19.5</points>
<intersection>54.5 1</intersection>
<intersection>60.5 8</intersection>
<intersection>76.5 10</intersection>
<intersection>100 12</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>54.5,-8,57,-8</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>54.5 1</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>60.5,-21,60.5,-19.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>76.5,-21,76.5,-19.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>100,-21,100,-19.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>17</ID>
<points>54.5,-62.5,142,-62.5</points>
<intersection>54.5 1</intersection>
<intersection>142 18</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>142,-62.5,142,-52</points>
<connection>
<GID>7</GID>
<name>N_in2</name></connection>
<intersection>-62.5 17</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>39,-21,116.5,-21</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>54.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-13.5,43.5,-12</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>-13.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>47.5,-21,47.5,-13.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>43.5,-13.5,112.5,-13.5</points>
<intersection>43.5 0</intersection>
<intersection>47.5 1</intersection>
<intersection>112.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>112.5,-21,112.5,-13.5</points>
<connection>
<GID>11</GID>
<name>IN_2</name></connection>
<intersection>-13.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-16,57,-12</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>-16 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>53,-21,53,-16</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-16,126.5,-16</points>
<intersection>31.5 13</intersection>
<intersection>53 1</intersection>
<intersection>57 0</intersection>
<intersection>69 4</intersection>
<intersection>90.5 6</intersection>
<intersection>109 11</intersection>
<intersection>126.5 9</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>69,-21,69,-16</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>-16 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>90.5,-21,90.5,-16</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-16 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>126.5,-38,126.5,-16</points>
<intersection>-38 10</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>126.5,-38,129,-38</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>126.5 9</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>109,-21,109,-16</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-16 2</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>31.5,-21,31.5,-16</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-16 2</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-21,56.5,-14.5</points>
<connection>
<GID>19</GID>
<name>IN_2</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>38.5,-14.5,38.5,-12</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-14.5,56.5,-14.5</points>
<intersection>38.5 1</intersection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-27.5,50,-27</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-27,50,-27</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-27.5,52,-27</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<connection>
<GID>18</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-27.5,54,-27</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54,-27,58.5,-27</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-27.5,70.5,-27</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>68,-27,70.5,-27</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-27.5,72.5,-27</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>72.5,-27,74.5,-27</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-58.5,45.5,-8</points>
<intersection>-58.5 9</intersection>
<intersection>-21 11</intersection>
<intersection>-17.5 2</intersection>
<intersection>-8 7</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>72.5,-21,72.5,-17.5</points>
<connection>
<GID>28</GID>
<name>IN_2</name></connection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-17.5,83,-17.5</points>
<intersection>45.5 0</intersection>
<intersection>72.5 1</intersection>
<intersection>83 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>83,-21,83,-17.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>45.5,-8,48,-8</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>45.5,-58.5,103,-58.5</points>
<intersection>45.5 0</intersection>
<intersection>103 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>103,-58.5,103,-51.5</points>
<connection>
<GID>5</GID>
<name>N_in2</name></connection>
<intersection>-58.5 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>45.5,-21,88.5,-21</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-60.5,50,-8</points>
<intersection>-60.5 13</intersection>
<intersection>-21 15</intersection>
<intersection>-19 2</intersection>
<intersection>-8 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>74.5,-21,74.5,-19</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>50,-19,98,-19</points>
<intersection>50 0</intersection>
<intersection>74.5 1</intersection>
<intersection>98 8</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50,-8,52.5,-8</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>98,-21,98,-19</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>50,-60.5,124.5,-60.5</points>
<intersection>50 0</intersection>
<intersection>124.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>124.5,-60.5,124.5,-52</points>
<connection>
<GID>9</GID>
<name>N_in2</name></connection>
<intersection>-60.5 13</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>50,-21,107,-21</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-15.5,52.5,-12</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>85,-21,85,-15.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>26,-15.5,114.5,-15.5</points>
<intersection>26 6</intersection>
<intersection>52.5 0</intersection>
<intersection>85 1</intersection>
<intersection>114.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>114.5,-21,114.5,-15.5</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>26,-21,26,-15.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-15.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-14,33.5,-12</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-14 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>94,-21,94,-14</points>
<connection>
<GID>32</GID>
<name>IN_3</name></connection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-14,94,-14</points>
<intersection>33.5 0</intersection>
<intersection>94 1</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-15,48,-12</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>96,-21,96,-15</points>
<connection>
<GID>32</GID>
<name>IN_2</name></connection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>48,-15,96,-15</points>
<intersection>48 0</intersection>
<intersection>96 1</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-27.5,89.5,-27</points>
<connection>
<GID>33</GID>
<name>IN_1</name></connection>
<connection>
<GID>31</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-27.5,91.5,-27</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-27,97,-27</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>91.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-27.5,87.5,-27</points>
<connection>
<GID>33</GID>
<name>IN_2</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>84,-27,87.5,-27</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>87.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-38,52,-33.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-38,54.5,-38</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-38,71.5,-33.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-38,74,-38</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-38,89.5,-33.5</points>
<connection>
<GID>33</GID>
<name>OUT</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-38,93,-38</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-35,129,-35</points>
<intersection>33.5 3</intersection>
<intersection>54.5 5</intersection>
<intersection>74 7</intersection>
<intersection>93 9</intersection>
<intersection>111 15</intersection>
<intersection>129 17</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33.5,-41,33.5,-35</points>
<intersection>-41 24</intersection>
<intersection>-35 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>54.5,-41,54.5,-35</points>
<connection>
<GID>35</GID>
<name>clock</name></connection>
<intersection>-35 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>74,-41,74,-35</points>
<connection>
<GID>36</GID>
<name>clock</name></connection>
<intersection>-35 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>93,-41,93,-35</points>
<connection>
<GID>37</GID>
<name>clock</name></connection>
<intersection>-35 1</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>111,-41,111,-35</points>
<connection>
<GID>8</GID>
<name>clock</name></connection>
<intersection>-35 1</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>129,-41,129,-35</points>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>30,-41,34.5,-41</points>
<connection>
<GID>34</GID>
<name>clock</name></connection>
<connection>
<GID>40</GID>
<name>CLK</name></connection>
<intersection>33.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-36,37.5,-34</points>
<connection>
<GID>34</GID>
<name>set</name></connection>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>-36 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>37.5,-36,96,-36</points>
<connection>
<GID>37</GID>
<name>set</name></connection>
<connection>
<GID>36</GID>
<name>set</name></connection>
<connection>
<GID>35</GID>
<name>set</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-45.5,37.5,-44</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-44,96,-44</points>
<connection>
<GID>37</GID>
<name>clear</name></connection>
<connection>
<GID>36</GID>
<name>clear</name></connection>
<connection>
<GID>35</GID>
<name>clear</name></connection>
<connection>
<GID>34</GID>
<name>clear</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-50,43.5,-38</points>
<connection>
<GID>2</GID>
<name>N_in3</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-38,43.5,-38</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-50,65,-38</points>
<connection>
<GID>3</GID>
<name>N_in3</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60.5,-38,65,-38</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-50,86,-38</points>
<connection>
<GID>4</GID>
<name>N_in3</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-38,86,-38</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-49.5,103,-38</points>
<connection>
<GID>5</GID>
<name>N_in3</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-38,103,-38</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-50,142,-38</points>
<connection>
<GID>7</GID>
<name>N_in3</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-38,142,-38</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-50,124.5,-38</points>
<connection>
<GID>9</GID>
<name>N_in3</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,-38,124.5,-38</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-27.5,110.5,-27</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>108,-27,110.5,-27</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-27.5,112.5,-27</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>112.5,-27,114.5,-27</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<intersection>112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-38,111.5,-33.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-38,111.5,-38</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-27.5,30.5,-27</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<connection>
<GID>14</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-27.5,28.5,-27</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>25,-27,28.5,-27</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-27.5,32.5,-27</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-27,37,-27</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-38,30.5,-33.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-38,34.5,-38</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 1>
<page 2>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 2>
<page 3>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 3>
<page 4>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 4>
<page 5>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 5>
<page 6>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 6>
<page 7>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 7>
<page 8>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 8>
<page 9>
<PageViewport>0,0,44.2,-46.1</PageViewport></page 9></circuit>