<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-150.586,31.6173,289.986,-189.933</PageViewport>
<gate>
<ID>1</ID>
<type>AE_SMALL_INVERTER</type>
<position>-74,-26</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>-78,-23.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3</ID>
<type>AE_SMALL_INVERTER</type>
<position>-74,-33.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-78,-31</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_DFF_LOW</type>
<position>-68,0.5</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>3 </output>
<input>
<ID>clear</ID>2 </input>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_SMALL_INVERTER</type>
<position>-62,-6.5</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_DFF_LOW</type>
<position>-68,-10</position>
<input>
<ID>IN_0</ID>19 </input>
<output>
<ID>OUT_0</ID>7 </output>
<input>
<ID>clear</ID>2 </input>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_AND2</type>
<position>-51,3.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>-87.5,-3</position>
<gparam>LABEL_TEXT Clock</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>-87,-13.5</position>
<gparam>LABEL_TEXT RST</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>-84,-23</position>
<gparam>LABEL_TEXT M1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>-51,-1</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_AND3</type>
<position>-51,-6.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>8 </input>
<input>
<ID>IN_2</ID>9 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>-84,-30.5</position>
<gparam>LABEL_TEXT M0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AE_SMALL_INVERTER</type>
<position>-62,4</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_OR3</type>
<position>-41.5,-1</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>12 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_AND4</type>
<position>-48,-16.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>8 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND3</type>
<position>-48,-24</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>9 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_AND3</type>
<position>-48,-30.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_AND4</type>
<position>-48,-38</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>14 </input>
<input>
<ID>IN_2</ID>8 </input>
<input>
<ID>IN_3</ID>9 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>21</ID>
<type>AE_OR4</type>
<position>-40.5,-27</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>17 </input>
<input>
<ID>IN_3</ID>18 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>-46,-46</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND3</type>
<position>-46,-51.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_OR2</type>
<position>-40,-48.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>GA_LED</type>
<position>-34.5,-48.5</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>-31,-48</position>
<gparam>LABEL_TEXT G</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_AND3</type>
<position>-44.5,-59.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>5 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>-34.5,-59.5</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>-31,-59</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>-82,-14</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_SMALL_INVERTER</type>
<position>-76,-13.5</position>
<input>
<ID>IN_0</ID>24 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-82,-3.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>-62.5,2</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>-62.5,-9</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-73.5,-11,-73.5,-0.5</points>
<intersection>-11 3</intersection>
<intersection>-3.5 4</intersection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-73.5,-0.5,-71,-0.5</points>
<connection>
<GID>5</GID>
<name>clock</name></connection>
<intersection>-73.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-73.5,-11,-71,-11</points>
<connection>
<GID>7</GID>
<name>clock</name></connection>
<intersection>-73.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-80,-3.5,-73.5,-3.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-72.5,-15,-72.5,-3.5</points>
<intersection>-15 1</intersection>
<intersection>-13.5 6</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72.5,-15,-68,-15</points>
<intersection>-72.5 0</intersection>
<intersection>-68 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-72.5,-3.5,-68,-3.5</points>
<connection>
<GID>5</GID>
<name>clear</name></connection>
<intersection>-72.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-68,-15,-68,-14</points>
<connection>
<GID>7</GID>
<name>clear</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-74,-13.5,-72.5,-13.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>-72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-64.5,-57.5,-64.5,4</points>
<intersection>-57.5 13</intersection>
<intersection>-49.5 11</intersection>
<intersection>-45 9</intersection>
<intersection>-35 7</intersection>
<intersection>-28.5 5</intersection>
<intersection>-4.5 3</intersection>
<intersection>2.5 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64.5,4,-64,4</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-65,2.5,-64.5,2.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-64.5,-4.5,-54,-4.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-64.5,-28.5,-51,-28.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-64.5,-35,-51,-35</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-64.5,-45,-49,-45</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-64.5,-49.5,-49,-49.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-64.5,-57.5,-47.5,-57.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>-64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57,-22,-57,4.5</points>
<intersection>-22 6</intersection>
<intersection>-13.5 4</intersection>
<intersection>4 1</intersection>
<intersection>4.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60,4,-57,4</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,4.5,-54,4.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-57,-13.5,-51,-13.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>-57 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-57,-22,-51,-22</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-57 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,-61.5,-57.5,2.5</points>
<intersection>-61.5 8</intersection>
<intersection>-47 6</intersection>
<intersection>-23.5 2</intersection>
<intersection>2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57.5,2.5,-54,2.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-76,-23.5,-57.5,-23.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>-76 4</intersection>
<intersection>-57.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-76,-26,-76,-23.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-57.5,-47,-49,-47</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-57.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-57.5,-61.5,-47.5,-61.5</points>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<intersection>-57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-56.5,-53.5,-56.5,-2</points>
<intersection>-53.5 8</intersection>
<intersection>-32.5 6</intersection>
<intersection>-31 2</intersection>
<intersection>-19.5 5</intersection>
<intersection>-2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56.5,-2,-54,-2</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>-56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-76,-31,-56.5,-31</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-76 4</intersection>
<intersection>-56.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-76,-33.5,-76,-31</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-56.5,-19.5,-51,-19.5</points>
<connection>
<GID>17</GID>
<name>IN_3</name></connection>
<intersection>-56.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-56.5,-32.5,-51,-32.5</points>
<connection>
<GID>19</GID>
<name>IN_2</name></connection>
<intersection>-56.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-56.5,-53.5,-49,-53.5</points>
<connection>
<GID>23</GID>
<name>IN_2</name></connection>
<intersection>-56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-65,-8,-58.5,-8</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-64 5</intersection>
<intersection>-58.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-58.5,-8,-58.5,0</points>
<intersection>-8 1</intersection>
<intersection>0 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-58.5,0,-54,0</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-58.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-64,-59.5,-64,-6.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-59.5 13</intersection>
<intersection>-51.5 11</intersection>
<intersection>-30.5 9</intersection>
<intersection>-24 7</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-64,-24,-51,-24</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>-64 5</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-64,-30.5,-51,-30.5</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>-64 5</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-64,-51.5,-49,-51.5</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>-64 5</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-64,-59.5,-47.5,-59.5</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>-64 5</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55.5,-39,-55.5,-6.5</points>
<intersection>-39 4</intersection>
<intersection>-26 1</intersection>
<intersection>-17.5 3</intersection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72,-26,-55.5,-26</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>-55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-55.5,-6.5,-54,-6.5</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>-55.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-55.5,-17.5,-51,-17.5</points>
<connection>
<GID>17</GID>
<name>IN_2</name></connection>
<intersection>-55.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-55.5,-39,-51,-39</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>-55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54.5,-41,-54.5,-8.5</points>
<intersection>-41 4</intersection>
<intersection>-33.5 1</intersection>
<intersection>-26 3</intersection>
<intersection>-8.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-72,-33.5,-54.5,-33.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-54.5,-8.5,-54,-8.5</points>
<connection>
<GID>13</GID>
<name>IN_2</name></connection>
<intersection>-54.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-54.5,-26,-51,-26</points>
<connection>
<GID>18</GID>
<name>IN_2</name></connection>
<intersection>-54.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-54.5,-41,-51,-41</points>
<connection>
<GID>20</GID>
<name>IN_3</name></connection>
<intersection>-54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48,-1,-44.5,-1</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<connection>
<GID>12</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,1,-46.5,3.5</points>
<intersection>1 1</intersection>
<intersection>3.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-46.5,1,-44.5,1</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-48,3.5,-46.5,3.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>-46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46.5,-6.5,-46.5,-3</points>
<intersection>-6.5 2</intersection>
<intersection>-3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-46.5,-3,-44.5,-3</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<intersection>-46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-48,-6.5,-46.5,-6.5</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>-46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-71,2.5,-71,10</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>10 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-71,10,-38.5,10</points>
<intersection>-71 0</intersection>
<intersection>-38.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-38.5,-1,-38.5,10</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>10 2</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-55.5,-15.5,-55.5,-6.5</points>
<intersection>-15.5 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60,-6.5,-55.5,-6.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-55.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-57,-15.5,-51,-15.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>-57 3</intersection>
<intersection>-55.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-57,-37,-57,-15.5</points>
<intersection>-37 4</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-57,-37,-51,-37</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-57 3</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43.5,-24,-43.5,-16.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-45,-16.5,-43.5,-16.5</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>-43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,-26,-44.5,-24</points>
<intersection>-26 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44.5,-26,-43.5,-26</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-45,-24,-44.5,-24</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,-30.5,-44.5,-28</points>
<intersection>-30.5 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44.5,-28,-43.5,-28</points>
<connection>
<GID>21</GID>
<name>IN_2</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-45,-30.5,-44.5,-30.5</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43.5,-38,-43.5,-30</points>
<connection>
<GID>21</GID>
<name>IN_3</name></connection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45,-38,-43.5,-38</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>-43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75,-8,-75,12</points>
<intersection>-8 1</intersection>
<intersection>12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-75,-8,-71,-8</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>-75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-75,12,-36.5,12</points>
<intersection>-75 0</intersection>
<intersection>-36.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-36.5,-27,-36.5,12</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>12 2</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-47.5,-43,-46</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<connection>
<GID>22</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-51.5,-43,-49.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<connection>
<GID>23</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-37,-48.5,-35.5,-48.5</points>
<connection>
<GID>25</GID>
<name>N_in0</name></connection>
<connection>
<GID>24</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41.5,-59.5,-35.5,-59.5</points>
<connection>
<GID>28</GID>
<name>N_in0</name></connection>
<connection>
<GID>27</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80,-14,-78,-14</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>-78 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-78,-14,-78,-13.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-14 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-95.5148,-0.0370359,234.915,-166.2</PageViewport></page 1>
<page 2>
<PageViewport>-23.2333,11.6667,162.633,-81.8</PageViewport></page 2>
<page 3>
<PageViewport>0,1.16081e-006,139.4,-70.1</PageViewport></page 3>
<page 4>
<PageViewport>0,1.16081e-006,139.4,-70.1</PageViewport></page 4>
<page 5>
<PageViewport>0,1.16081e-006,139.4,-70.1</PageViewport></page 5>
<page 6>
<PageViewport>0,1.16081e-006,139.4,-70.1</PageViewport></page 6>
<page 7>
<PageViewport>0,1.16081e-006,139.4,-70.1</PageViewport></page 7>
<page 8>
<PageViewport>0,1.16081e-006,139.4,-70.1</PageViewport></page 8>
<page 9>
<PageViewport>0,1.16081e-006,139.4,-70.1</PageViewport></page 9></circuit>