<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-36.2605,-1.06592,102.71,-70.9501</PageViewport>
<gate>
<ID>1</ID>
<type>BB_CLOCK</type>
<position>21.5,-20</position>
<output>
<ID>CLK</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>2</ID>
<type>DE_TO</type>
<position>29,-20</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>21.5,-25.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>DE_TO</type>
<position>29,-25</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /MR0</lparam></gate>
<gate>
<ID>5</ID>
<type>DE_TO</type>
<position>29,-27.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /MR1</lparam></gate>
<gate>
<ID>6</ID>
<type>DE_TO</type>
<position>29,-30</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /MR2</lparam></gate>
<gate>
<ID>7</ID>
<type>DE_TO</type>
<position>29,-32.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /MR3</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>22.5,-38.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>DE_TO</type>
<position>29,-39</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Load</lparam></gate>
<gate>
<ID>10</ID>
<type>DE_TO</type>
<position>29,-43</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>22,-43</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>27.5,-56</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>8 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>13</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>46,-56</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>10 </input>
<input>
<ID>IN_3</ID>9 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>14</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>64,-56</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>15 </input>
<input>
<ID>IN_2</ID>14 </input>
<input>
<ID>IN_3</ID>13 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>15</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>82.5,-56</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>18 </input>
<input>
<ID>IN_3</ID>17 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 4</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>19,-52.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q3_3</lparam></gate>
<gate>
<ID>17</ID>
<type>DA_FROM</type>
<position>19,-55</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q3_2</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>19,-57.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q3_1</lparam></gate>
<gate>
<ID>19</ID>
<type>DA_FROM</type>
<position>19,-60</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q3_0</lparam></gate>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>36,-52.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q2_3</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>36,-55</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q2_2</lparam></gate>
<gate>
<ID>22</ID>
<type>DA_FROM</type>
<position>36,-57.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q2_1</lparam></gate>
<gate>
<ID>23</ID>
<type>DA_FROM</type>
<position>36,-60</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q2_0</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>54.5,-52.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q1_3</lparam></gate>
<gate>
<ID>25</ID>
<type>DA_FROM</type>
<position>54.5,-55</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q1_2</lparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>54.5,-57.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q1_1</lparam></gate>
<gate>
<ID>27</ID>
<type>DA_FROM</type>
<position>54.5,-60</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q1_0</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>73,-52.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q0_3</lparam></gate>
<gate>
<ID>29</ID>
<type>DA_FROM</type>
<position>73,-55</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q0_2</lparam></gate>
<gate>
<ID>30</ID>
<type>DA_FROM</type>
<position>73,-57.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q0_1</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>73,-60</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q0_0</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>14.5,-19.5</position>
<gparam>LABEL_TEXT Clock</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>15,-25</position>
<gparam>LABEL_TEXT /Reset</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>16.5,-38</position>
<gparam>LABEL_TEXT /Load</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>17,-42.5</position>
<gparam>LABEL_TEXT CE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>21,-3.5</position>
<gparam>LABEL_TEXT Minute : Page2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>22.5,-7.5</position>
<gparam>LABEL_TEXT Hour : Page3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-20,27,-20</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>1</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23.5,-25.5,27,-25.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>27 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27,-32.5,27,-25</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-25.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-38.5,27,-38.5</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>27 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>27,-39,27,-38.5</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>-38.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-43,27,-43</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-60,22.5,-57</points>
<intersection>-60 2</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-57,24.5,-57</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-60,22.5,-60</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-57.5,22.5,-56</points>
<intersection>-57.5 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-56,24.5,-56</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-57.5,22.5,-57.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-55,24.5,-55</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-54,22.5,-52.5</points>
<intersection>-54 1</intersection>
<intersection>-52.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-54,24.5,-54</points>
<connection>
<GID>12</GID>
<name>IN_3</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-52.5,22.5,-52.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-54,40.5,-52.5</points>
<intersection>-54 1</intersection>
<intersection>-52.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-54,43,-54</points>
<connection>
<GID>13</GID>
<name>IN_3</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-52.5,40.5,-52.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-55,43,-55</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-57.5,40.5,-56</points>
<intersection>-57.5 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-56,43,-56</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-57.5,40.5,-57.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-60,40.5,-57</points>
<intersection>-60 2</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-57,43,-57</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-60,40.5,-60</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-54,58.5,-52.5</points>
<intersection>-54 1</intersection>
<intersection>-52.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-54,61,-54</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-52.5,58.5,-52.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,-55,61,-55</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-57.5,58.5,-56</points>
<intersection>-57.5 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-56,61,-56</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-57.5,58.5,-57.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-60,58.5,-57</points>
<intersection>-60 2</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-57,61,-57</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-60,58.5,-60</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-54,77,-52.5</points>
<intersection>-54 1</intersection>
<intersection>-52.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-54,79.5,-54</points>
<connection>
<GID>15</GID>
<name>IN_3</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-52.5,77,-52.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-55,79.5,-55</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<connection>
<GID>15</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-57.5,77,-56</points>
<intersection>-57.5 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-56,79.5,-56</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-57.5,77,-57.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-60,77,-57</points>
<intersection>-60 2</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-57,79.5,-57</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-60,77,-60</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-27.7986,75.4025,407.243,-143.367</PageViewport>
<gate>
<ID>194</ID>
<type>AE_OR2</type>
<position>134,10</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>161 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>198</ID>
<type>AE_OR2</type>
<position>78,-2.5</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>163 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AF_DFF_LOW</type>
<position>9.5,-16.5</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUTINV_0</ID>25 </output>
<output>
<ID>OUT_0</ID>21 </output>
<input>
<ID>clear</ID>157 </input>
<input>
<ID>clock</ID>69 </input>
<input>
<ID>clock_enable</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>37</ID>
<type>AF_DFF_LOW</type>
<position>24,-16.5</position>
<input>
<ID>IN_0</ID>84 </input>
<output>
<ID>OUTINV_0</ID>26 </output>
<output>
<ID>OUT_0</ID>23 </output>
<input>
<ID>clear</ID>157 </input>
<input>
<ID>clock</ID>69 </input>
<input>
<ID>clock_enable</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>38</ID>
<type>AF_DFF_LOW</type>
<position>38,-16.5</position>
<input>
<ID>IN_0</ID>82 </input>
<output>
<ID>OUTINV_0</ID>22 </output>
<output>
<ID>OUT_0</ID>24 </output>
<input>
<ID>clear</ID>157 </input>
<input>
<ID>clock</ID>69 </input>
<input>
<ID>clock_enable</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_AND2</type>
<position>9,-35.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND2</type>
<position>14,-35.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_AND2</type>
<position>23.5,-35.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_AND3</type>
<position>29.5,-35.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>26 </input>
<input>
<ID>IN_2</ID>25 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>43</ID>
<type>AE_OR2</type>
<position>11.5,-42</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AE_OR2</type>
<position>26.5,-42</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>16.5,20.5</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q1_2</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>29,20</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q1_1</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>42.5,20</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q1_0</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>4.5,20</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q1_3</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>-1.5,20</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>AF_DFF_LOW</type>
<position>84.5,-23.5</position>
<input>
<ID>IN_0</ID>158 </input>
<output>
<ID>OUTINV_0</ID>41 </output>
<output>
<ID>OUT_0</ID>34 </output>
<input>
<ID>clear</ID>156 </input>
<input>
<ID>clock</ID>52 </input>
<input>
<ID>clock_enable</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>51</ID>
<type>AF_DFF_LOW</type>
<position>99,-23.5</position>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUTINV_0</ID>40 </output>
<output>
<ID>OUT_0</ID>37 </output>
<input>
<ID>clear</ID>156 </input>
<input>
<ID>clock</ID>52 </input>
<input>
<ID>clock_enable</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>52</ID>
<type>AF_DFF_LOW</type>
<position>113,-23.5</position>
<input>
<ID>IN_0</ID>160 </input>
<output>
<ID>OUTINV_0</ID>35 </output>
<output>
<ID>OUT_0</ID>38 </output>
<input>
<ID>clear</ID>156 </input>
<input>
<ID>clock</ID>52 </input>
<input>
<ID>clock_enable</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>53</ID>
<type>AF_DFF_LOW</type>
<position>128,-23.5</position>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUTINV_0</ID>99 </output>
<output>
<ID>OUT_0</ID>39 </output>
<input>
<ID>clear</ID>156 </input>
<input>
<ID>clock</ID>52 </input>
<input>
<ID>clock_enable</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_AND3</type>
<position>93.5,-43</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>37 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_AND3</type>
<position>87,-43</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>35 </input>
<input>
<ID>IN_2</ID>34 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_AND3</type>
<position>104,-43</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>40 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_LABEL</type>
<position>93.5,34.5</position>
<gparam>LABEL_TEXT Q0_3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_AND3</type>
<position>110.5,-43</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>41 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_LABEL</type>
<position>107,34</position>
<gparam>LABEL_TEXT Q0_2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_AND3</type>
<position>117,-43</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>41 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_LABEL</type>
<position>122.5,34</position>
<gparam>LABEL_TEXT Q0_1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_AND3</type>
<position>127.5,-43</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>35 </input>
<input>
<ID>IN_2</ID>41 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_LABEL</type>
<position>136.5,33</position>
<gparam>LABEL_TEXT Q0_0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_AND2</type>
<position>133,-43</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_LABEL</type>
<position>42.5,46</position>
<gparam>LABEL_TEXT Q1_0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AE_OR2</type>
<position>90.5,-50</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>151 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_LABEL</type>
<position>28,46</position>
<gparam>LABEL_TEXT Q1_1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AE_OR3</type>
<position>110.5,-50</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>44 </input>
<input>
<ID>IN_2</ID>45 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>256</ID>
<type>AA_LABEL</type>
<position>14.5,45.5</position>
<gparam>LABEL_TEXT Q1_2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AE_OR2</type>
<position>130.5,-49.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>68.5,-23.5</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>65</ID>
<type>DE_TO</type>
<position>91.5,0</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q0_3</lparam></gate>
<gate>
<ID>66</ID>
<type>DE_TO</type>
<position>106,0</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q0_2</lparam></gate>
<gate>
<ID>67</ID>
<type>DE_TO</type>
<position>119,0</position>
<input>
<ID>IN_0</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q0_1</lparam></gate>
<gate>
<ID>68</ID>
<type>DE_TO</type>
<position>133,0</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q0_0</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND2</type>
<position>-41.5,-67</position>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>BM_NORX4</type>
<position>-60,-48</position>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_AND2</type>
<position>35.5,29.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_AND2</type>
<position>51,-68.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>93,27.5</position>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_AND2</type>
<position>71.5,-68</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>BM_NORX3</type>
<position>-26.5,-60</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_AND2</type>
<position>59.5,-78.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AE_SMALL_INVERTER</type>
<position>69.5,32.5</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>13,40.5</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>28,40.5</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>85</ID>
<type>AE_SMALL_INVERTER</type>
<position>91,25</position>
<input>
<ID>IN_0</ID>126 </input>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>86</ID>
<type>BE_NOR2</type>
<position>-49,-25</position>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>87</ID>
<type>AA_TOGGLE</type>
<position>42,41</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>88</ID>
<type>DA_FROM</type>
<position>44.5,-82.5</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /MR1</lparam></gate>
<gate>
<ID>90</ID>
<type>DA_FROM</type>
<position>71.5,-56.5</position>
<input>
<ID>IN_0</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /MR0</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_SMALL_INVERTER</type>
<position>11,38.5</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>66 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>92</ID>
<type>DA_FROM</type>
<position>-12,9.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>94</ID>
<type>DA_FROM</type>
<position>69,3</position>
<input>
<ID>IN_0</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>95</ID>
<type>AE_SMALL_INVERTER</type>
<position>26,39</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>96</ID>
<type>AE_OR2</type>
<position>8.5,27</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_SMALL_INVERTER</type>
<position>39.5,39</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>98</ID>
<type>DA_FROM</type>
<position>-6.5,-16.5</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>100</ID>
<type>DA_FROM</type>
<position>-13,55.5</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID /Load</lparam></gate>
<gate>
<ID>102</ID>
<type>AE_SMALL_INVERTER</type>
<position>-24.5,-52.5</position>
<gparam>angle 0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_AND2</type>
<position>4,33</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_AND2</type>
<position>-1,7</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AE_OR2</type>
<position>25.5,24.5</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>AE_OR2</type>
<position>38.5,24.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_AND2</type>
<position>21.5,30.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_AND2</type>
<position>-46,-66</position>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_AND2</type>
<position>27,32.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>114</ID>
<type>AA_AND2</type>
<position>-7,49</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_AND2</type>
<position>12,33</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_AND2</type>
<position>41,32.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_SMALL_INVERTER</type>
<position>-13,2.5</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_AND2</type>
<position>92,19.5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>AE_OR2</type>
<position>1,1.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND2</type>
<position>130.5,16</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_TOGGLE</type>
<position>108,27</position>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>152</ID>
<type>DE_TO</type>
<position>70.5,-83</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID H_change</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_TOGGLE</type>
<position>123,27</position>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_TOGGLE</type>
<position>137,27.5</position>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>156</ID>
<type>AE_SMALL_INVERTER</type>
<position>106,25</position>
<input>
<ID>IN_0</ID>126 </input>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>157</ID>
<type>AE_SMALL_INVERTER</type>
<position>121,25.5</position>
<input>
<ID>IN_0</ID>126 </input>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>159</ID>
<type>AE_OR2</type>
<position>103.5,13.5</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>AE_SMALL_INVERTER</type>
<position>134.5,25.5</position>
<input>
<ID>IN_0</ID>126 </input>
<output>
<ID>OUT_0</ID>121 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>163</ID>
<type>DA_FROM</type>
<position>67.5,42</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID /Load</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_AND2</type>
<position>99,19.5</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_AND2</type>
<position>116.5,17</position>
<input>
<ID>IN_0</ID>147 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>142 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_AND2</type>
<position>123,18</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>AA_AND2</type>
<position>88,35.5</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>126 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_AND2</type>
<position>107,19.5</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>128 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_AND2</type>
<position>136,19</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_AND2</type>
<position>86,19</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>184</ID>
<type>AE_OR2</type>
<position>89.5,12</position>
<input>
<ID>IN_0</ID>136 </input>
<input>
<ID>IN_1</ID>135 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>AE_OR2</type>
<position>121,10.5</position>
<input>
<ID>IN_0</ID>141 </input>
<input>
<ID>IN_1</ID>142 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-23,14,20.5</points>
<intersection>-23 2</intersection>
<intersection>-14.5 1</intersection>
<intersection>20.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12.5,-14.5,14,-14.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-23,14,-23</points>
<intersection>8 3</intersection>
<intersection>14 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>8,-69.5,8,-23</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>-69.5 5</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>14,20.5,14.5,20.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>8,-69.5,48,-69.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>8 3</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-32.5,10,-30</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-30,41,-30</points>
<intersection>10 0</intersection>
<intersection>24.5 4</intersection>
<intersection>41 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>41,-45,41,-17.5</points>
<connection>
<GID>38</GID>
<name>OUTINV_0</name></connection>
<intersection>-45 19</intersection>
<intersection>-30 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>24.5,-32.5,24.5,-30</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>31.5,-45,41,-45</points>
<intersection>31.5 23</intersection>
<intersection>41 2</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>31.5,-45,31.5,31</points>
<intersection>-45 19</intersection>
<intersection>31 28</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>31.5,31,36.5,31</points>
<intersection>31.5 23</intersection>
<intersection>36.5 32</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>36.5,31,36.5,32.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>31 28</intersection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-24.5,28.5,-14.5</points>
<intersection>-24.5 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-14.5,28.5,-14.5</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>27 5</intersection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-24.5,28.5,-24.5</points>
<intersection>13 3</intersection>
<intersection>22.5 4</intersection>
<intersection>28.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13,-32.5,13,-24.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>-24.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>22.5,-32.5,22.5,-24.5</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>-24.5 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>27,-14.5,27,20</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>-14.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-32.5,15,-26</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-26,42.5,-26</points>
<intersection>15 0</intersection>
<intersection>31.5 4</intersection>
<intersection>42.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>42.5,-26,42.5,-14.5</points>
<intersection>-26 1</intersection>
<intersection>-14.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>40.5,-14.5,42.5,-14.5</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>40.5 5</intersection>
<intersection>42.5 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>31.5,-67.5,31.5,-26</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-67.5 6</intersection>
<intersection>-26 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>40.5,-14.5,40.5,20</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>-14.5 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>31.5,-67.5,48,-67.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>31.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-32.5,27.5,-27.5</points>
<connection>
<GID>42</GID>
<name>IN_2</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12.5,-27.5,27.5,-27.5</points>
<intersection>12.5 2</intersection>
<intersection>27.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>12.5,-27.5,12.5,-17.5</points>
<connection>
<GID>36</GID>
<name>OUTINV_0</name></connection>
<intersection>-27.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-32.5,29.5,-17.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-17.5,29.5,-17.5</points>
<connection>
<GID>37</GID>
<name>OUTINV_0</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-39,10.5,-38.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>9,-38.5,10.5,-38.5</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-39,12.5,-38.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-38.5,14,-38.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-39,25.5,-38.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-38.5,25.5,-38.5</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-39,27.5,-38.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-38.5,29.5,-38.5</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-75.5,58.5,-68.5</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-68.5,58.5,-68.5</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0.5,20,2.5,20</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-29.5,88.5,-21.5</points>
<intersection>-29.5 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-21.5,88.5,-21.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>86.5 4</intersection>
<intersection>88.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>85,-29.5,88.5,-29.5</points>
<intersection>85 3</intersection>
<intersection>88.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>85,-67,85,-29.5</points>
<connection>
<GID>55</GID>
<name>IN_2</name></connection>
<intersection>-67 6</intersection>
<intersection>-29.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>86.5,-21.5,86.5,0</points>
<intersection>-21.5 1</intersection>
<intersection>0 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>86.5,0,89.5,0</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>86.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>74.5,-67,85,-67</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<intersection>85 3</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-40,87,-37.5</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-37.5,127.5,-37.5</points>
<intersection>87 0</intersection>
<intersection>112.5 3</intersection>
<intersection>116 2</intersection>
<intersection>127.5 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>116,-37.5,116,-24.5</points>
<connection>
<GID>52</GID>
<name>OUTINV_0</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>112.5,-40,112.5,-37.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>127.5,-40,127.5,-37.5</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>-37.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-31,103,0</points>
<intersection>-31 2</intersection>
<intersection>-21.5 1</intersection>
<intersection>0 9</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-21.5,103,-21.5</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-31,117,-31</points>
<intersection>91.5 3</intersection>
<intersection>103 0</intersection>
<intersection>110.5 6</intersection>
<intersection>117 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>91.5,-40,91.5,-31</points>
<connection>
<GID>54</GID>
<name>IN_2</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>110.5,-40,110.5,-31</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>117,-40,117,-31</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>-31 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>103,0,104,0</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-32,117.5,-21.5</points>
<intersection>-32 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-21.5,117.5,-21.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>115.5 7</intersection>
<intersection>117.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,-32,132,-32</points>
<intersection>93.5 3</intersection>
<intersection>104 4</intersection>
<intersection>117.5 0</intersection>
<intersection>132 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>93.5,-40,93.5,-32</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>104,-40,104,-32</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>132,-40,132,-32</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>115.5,-21.5,115.5,0</points>
<intersection>-21.5 1</intersection>
<intersection>0 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>115.5,0,117,0</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>115.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-33,131,0</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-33,131,-33</points>
<intersection>95.5 3</intersection>
<intersection>106 4</intersection>
<intersection>129.5 5</intersection>
<intersection>131 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>95.5,-69,95.5,-33</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>-69 6</intersection>
<intersection>-33 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>106,-40,106,-33</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>-33 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>129.5,-40,129.5,-33</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>74.5,-69,95.5,-69</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>95.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-40,102,-24.5</points>
<connection>
<GID>51</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>56</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-40,108.5,-35.5</points>
<connection>
<GID>57</GID>
<name>IN_2</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87.5,-35.5,125.5,-35.5</points>
<intersection>87.5 2</intersection>
<intersection>108.5 0</intersection>
<intersection>115 4</intersection>
<intersection>125.5 6</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>87.5,-35.5,87.5,-24.5</points>
<connection>
<GID>50</GID>
<name>OUTINV_0</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>115,-40,115,-35.5</points>
<connection>
<GID>58</GID>
<name>IN_2</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>125.5,-40,125.5,-35.5</points>
<connection>
<GID>59</GID>
<name>IN_2</name></connection>
<intersection>-35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91.5,-47,91.5,-46.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>93.5,-46.5,93.5,-46</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>91.5,-46.5,93.5,-46.5</points>
<intersection>91.5 0</intersection>
<intersection>93.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-47,89.5,-46.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>87,-46.5,87,-46</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>87,-46.5,89.5,-46.5</points>
<intersection>87 1</intersection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-47,110.5,-46</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<connection>
<GID>57</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-46.5,104,-46</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>108.5,-47,108.5,-46.5</points>
<connection>
<GID>62</GID>
<name>IN_2</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>104,-46.5,108.5,-46.5</points>
<intersection>104 0</intersection>
<intersection>108.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,-46.5,117,-46</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>112.5,-47,112.5,-46.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>112.5,-46.5,117,-46.5</points>
<intersection>112.5 1</intersection>
<intersection>117 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-46.5,129.5,-46</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-46,129.5,-46</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131.5,-46.5,131.5,-46</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>131.5,-46,133,-46</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>131.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-11,123.5,-11</points>
<intersection>70.5 10</intersection>
<intersection>80.5 9</intersection>
<intersection>92.5 8</intersection>
<intersection>109 7</intersection>
<intersection>123.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>123.5,-23.5,123.5,-11</points>
<intersection>-23.5 17</intersection>
<intersection>-11 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>109,-23.5,109,-11</points>
<intersection>-23.5 12</intersection>
<intersection>-11 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>92.5,-23.5,92.5,-11</points>
<intersection>-23.5 11</intersection>
<intersection>-11 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>80.5,-23.5,80.5,-11</points>
<intersection>-23.5 16</intersection>
<intersection>-11 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>70.5,-23.5,70.5,-11</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>92.5,-23.5,96,-23.5</points>
<connection>
<GID>51</GID>
<name>clock</name></connection>
<intersection>92.5 8</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>109,-23.5,110,-23.5</points>
<connection>
<GID>52</GID>
<name>clock</name></connection>
<intersection>109 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>80.5,-23.5,81.5,-23.5</points>
<connection>
<GID>50</GID>
<name>clock</name></connection>
<intersection>80.5 9</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>123.5,-23.5,125,-23.5</points>
<connection>
<GID>53</GID>
<name>clock</name></connection>
<intersection>123.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,35.5,42,39</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>60.5,-75.5,60.5,12.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>-68 14</intersection>
<intersection>12.5 11</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>-4,12.5,60.5,12.5</points>
<intersection>-4 12</intersection>
<intersection>60.5 6</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-4,8,-4,12.5</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>12.5 11</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>60.5,-68,68.5,-68</points>
<connection>
<GID>75</GID>
<name>OUT</name></connection>
<intersection>60.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,35.5,28,38.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,36,13,38.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,22.5,93,25.5</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<connection>
<GID>120</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>91,22.5,91,23</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<connection>
<GID>120</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,35.5,40,36</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>36 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>39.5,36,39.5,37</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>36 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>39.5,36,40,36</points>
<intersection>39.5 1</intersection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>26,35.5,26,37</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,36,11,36.5</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-7,43,-7,46</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>43 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-7,43,39.5,43</points>
<intersection>-7 1</intersection>
<intersection>11 4</intersection>
<intersection>26 6</intersection>
<intersection>39.5 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>11,40.5,11,43</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>43 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>26,41,26,43</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>43 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>39.5,41,39.5,43</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>43 2</intersection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27.5,2.5,-27.5,53</points>
<intersection>2.5 3</intersection>
<intersection>53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27.5,53,-8,53</points>
<intersection>-27.5 0</intersection>
<intersection>-11 5</intersection>
<intersection>-8 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-27.5,2.5,-15,2.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-27.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-11,53,-11,55.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>53 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-8,52,-8,53</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>53 1</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-4.5,-9,34,-9</points>
<intersection>-4.5 8</intersection>
<intersection>6 7</intersection>
<intersection>20.5 6</intersection>
<intersection>34 10</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>20.5,-16.5,20.5,-9</points>
<intersection>-16.5 13</intersection>
<intersection>-9 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>6,-16.5,6,-9</points>
<intersection>-16.5 12</intersection>
<intersection>-9 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-4.5,-16.5,-4.5,-9</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>-9 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>34,-16.5,34,-9</points>
<intersection>-16.5 11</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>34,-16.5,35,-16.5</points>
<connection>
<GID>38</GID>
<name>clock</name></connection>
<intersection>34 10</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>6,-16.5,6.5,-16.5</points>
<connection>
<GID>36</GID>
<name>clock</name></connection>
<intersection>6 7</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>20.5,-16.5,21,-16.5</points>
<connection>
<GID>37</GID>
<name>clock</name></connection>
<intersection>20.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6.5,-47.5,-6.5,39</points>
<intersection>-47.5 2</intersection>
<intersection>39 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>11.5,-47.5,11.5,-45</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>-47.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-6.5,-47.5,11.5,-47.5</points>
<intersection>-6.5 0</intersection>
<intersection>11.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-6.5,39,5,39</points>
<intersection>-6.5 0</intersection>
<intersection>5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>5,36,5,39</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>39 3</intersection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-6.5,22.5,33.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-6.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>26.5,-45,26.5,-6.5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>-6.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-6.5,26.5,-6.5</points>
<intersection>22.5 0</intersection>
<intersection>26.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9.5,30,12,30</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<connection>
<GID>96</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18.5,6,-4,6</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<intersection>-18.5 2</intersection>
<intersection>-4.5 10</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-18.5,6,-18.5,52</points>
<intersection>6 1</intersection>
<intersection>37 4</intersection>
<intersection>52 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-18.5,52,-6,52</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-18.5 2</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-18.5,37,3,37</points>
<intersection>-18.5 2</intersection>
<intersection>3 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>3,34.5,3,37</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>34.5 6</intersection>
<intersection>37 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>3,34.5,34.5,34.5</points>
<intersection>3 5</intersection>
<intersection>20.5 8</intersection>
<intersection>34.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>34.5,32.5,34.5,34.5</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>34.5 6</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>20.5,33.5,20.5,34.5</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>34.5 6</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-4.5,6,-4.5,9.5</points>
<intersection>6 1</intersection>
<intersection>9.5 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-10,9.5,-4.5,9.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>-4.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,30,7.5,30</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<connection>
<GID>96</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,7,32,7</points>
<intersection>5.5 5</intersection>
<intersection>19 4</intersection>
<intersection>32 7</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>19,-18.5,19,7</points>
<intersection>-18.5 9</intersection>
<intersection>7 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>5.5,-18.5,5.5,7</points>
<intersection>-18.5 10</intersection>
<intersection>1.5 11</intersection>
<intersection>7 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>32,-18.5,32,7</points>
<intersection>-18.5 8</intersection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>32,-18.5,35,-18.5</points>
<connection>
<GID>38</GID>
<name>clock_enable</name></connection>
<intersection>32 7</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>19,-18.5,21,-18.5</points>
<connection>
<GID>37</GID>
<name>clock_enable</name></connection>
<intersection>19 4</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>5.5,-18.5,6.5,-18.5</points>
<connection>
<GID>36</GID>
<name>clock_enable</name></connection>
<intersection>5.5 5</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>4,1.5,5.5,1.5</points>
<connection>
<GID>147</GID>
<name>OUT</name></connection>
<intersection>5.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21.5,27.5,24.5,27.5</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<connection>
<GID>106</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,28.5,27,29.5</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>28.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>26.5,27.5,26.5,28.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>28.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>26.5,28.5,27,28.5</points>
<intersection>26.5 1</intersection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,28.5,41,29.5</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>28.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>39.5,27.5,39.5,28.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>28.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>39.5,28.5,41,28.5</points>
<intersection>39.5 1</intersection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,26.5,35.5,27</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>27 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>37.5,27,37.5,27.5</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>27 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35.5,27,37.5,27</points>
<intersection>35.5 0</intersection>
<intersection>37.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-14.5,38.5,21.5</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-14.5,38.5,-14.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>59.5,-83,59.5,-81.5</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59.5,-83,68.5,-83</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>59.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-14.5,25.5,21.5</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-14.5,25.5,-14.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-14.5,8.5,24</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-14.5,8.5,-14.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,0.5,-7,2.5</points>
<intersection>0.5 1</intersection>
<intersection>2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7,0.5,-2,0.5</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>-7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-11,2.5,-7,2.5</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>-7 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,2.5,0,7</points>
<intersection>2.5 1</intersection>
<intersection>7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2,2.5,0,2.5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>0 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0,7,2,7</points>
<connection>
<GID>104</GID>
<name>OUT</name></connection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137,22,137,25.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>7</ID>
<points>89,-39,157.5,-39</points>
<intersection>89 35</intersection>
<intersection>119 9</intersection>
<intersection>134 10</intersection>
<intersection>157.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>157.5,-39,157.5,-24.5</points>
<intersection>-39 7</intersection>
<intersection>-24.5 32</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>119,-40,119,-39</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-39 7</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>134,-40,134,-39</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>-39 7</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>131,-24.5,157.5,-24.5</points>
<connection>
<GID>53</GID>
<name>OUTINV_0</name></connection>
<intersection>131.5 36</intersection>
<intersection>157.5 8</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>89,-40,89,-39</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>-39 7</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>131.5,-24.5,131.5,19</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>-24.5 32</intersection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,21,124,25</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>25 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>123,25,124,25</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>124 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,22.5,108,25</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<connection>
<GID>151</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,22,135,22.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>22.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>134.5,22.5,134.5,23.5</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>22.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>134.5,22.5,135,22.5</points>
<intersection>134.5 1</intersection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>122,21,122,23.5</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<intersection>23.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>121,23.5,122,23.5</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>122 6</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,22.5,106,23</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>88,29.5,88,32.5</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<intersection>29.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>88,29.5,134.5,29.5</points>
<intersection>88 1</intersection>
<intersection>91 10</intersection>
<intersection>106 4</intersection>
<intersection>121 6</intersection>
<intersection>134.5 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>106,27,106,29.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>29.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>121,27.5,121,29.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>29.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>134.5,27.5,134.5,29.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>29.5 2</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>91,27,91,29.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>29.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,39.5,87,39.5</points>
<intersection>84 5</intersection>
<intersection>87 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>84,39.5,84,42</points>
<intersection>39.5 1</intersection>
<intersection>42 8</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>87,38.5,87,39.5</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>39.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>67.5,42,84,42</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>67.5 9</intersection>
<intersection>84 5</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>67.5,32.5,67.5,42</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>42 8</intersection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,16.5,107,16.5</points>
<connection>
<GID>173</GID>
<name>OUT</name></connection>
<connection>
<GID>159</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>76.5,32,76.5,38.5</points>
<intersection>32 4</intersection>
<intersection>33.5 10</intersection>
<intersection>38.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>76.5,38.5,89,38.5</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>76.5 2</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>76.5,32,129.5,32</points>
<intersection>76.5 2</intersection>
<intersection>85 9</intersection>
<intersection>98 5</intersection>
<intersection>115.5 8</intersection>
<intersection>129.5 7</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>98,22.5,98,32</points>
<connection>
<GID>165</GID>
<name>IN_1</name></connection>
<intersection>32 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>129.5,19,129.5,32</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>32 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>115.5,20,115.5,32</points>
<connection>
<GID>167</GID>
<name>IN_1</name></connection>
<intersection>32 4</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>85,22,85,32</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<intersection>32 4</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>75.5,33.5,76.5,33.5</points>
<intersection>75.5 15</intersection>
<intersection>76.5 2</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>75.5,3,75.5,33.5</points>
<intersection>3 24</intersection>
<intersection>33.5 10</intersection></vsegment>
<hsegment>
<ID>24</ID>
<points>71,3,75.5,3</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>75 25</intersection>
<intersection>75.5 15</intersection></hsegment>
<vsegment>
<ID>25</ID>
<points>75,-3.5,75,3</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>3 24</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99,16.5,102.5,16.5</points>
<connection>
<GID>165</GID>
<name>OUT</name></connection>
<connection>
<GID>159</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,15,88.5,15.5</points>
<connection>
<GID>184</GID>
<name>IN_1</name></connection>
<intersection>15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>86,15.5,86,16</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<intersection>15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>86,15.5,88.5,15.5</points>
<intersection>86 1</intersection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,15.5,92,16.5</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<intersection>15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>90.5,15,90.5,15.5</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>90.5,15.5,92,15.5</points>
<intersection>90.5 1</intersection>
<intersection>92 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>130.5,13,133,13</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<connection>
<GID>194</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,14.5,136,16</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<intersection>14.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>135,13,135,14.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>14.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>135,14.5,136,14.5</points>
<intersection>135 1</intersection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,14,123,15</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<intersection>14 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>122,13.5,122,14</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>122,14,123,14</points>
<intersection>122 1</intersection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,13.5,116.5,14</points>
<connection>
<GID>167</GID>
<name>OUT</name></connection>
<intersection>13.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>116.5,13.5,120,13.5</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>130.5,-52.5,130.5,-16</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<intersection>-16 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>117.5,-16,117.5,20</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>117.5,-16,130.5,-16</points>
<intersection>117.5 1</intersection>
<intersection>130.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-53,106,-15</points>
<intersection>-53 4</intersection>
<intersection>-15 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>100,-15,100,22.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>100,-15,106,-15</points>
<intersection>100 1</intersection>
<intersection>106 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>106,-53,110.5,-53</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-53,90.5,-15.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>87,-15.5,87,22</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>87,-15.5,90.5,-15.5</points>
<intersection>87 1</intersection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-58,84.5,-27.5</points>
<connection>
<GID>50</GID>
<name>clear</name></connection>
<intersection>-58 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-58,84.5,-58</points>
<intersection>73.5 4</intersection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84.5,-27.5,128,-27.5</points>
<connection>
<GID>53</GID>
<name>clear</name></connection>
<connection>
<GID>52</GID>
<name>clear</name></connection>
<connection>
<GID>51</GID>
<name>clear</name></connection>
<intersection>84.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>73.5,-58,73.5,-56.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>-58 1</intersection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-4,-20.5,38,-20.5</points>
<connection>
<GID>38</GID>
<name>clear</name></connection>
<connection>
<GID>37</GID>
<name>clear</name></connection>
<connection>
<GID>36</GID>
<name>clear</name></connection>
<intersection>-4 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-4,-89,-4,-20.5</points>
<intersection>-89 6</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-4,-89,46.5,-89</points>
<intersection>-4 5</intersection>
<intersection>46.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>46.5,-89,46.5,-82.5</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>-89 6</intersection></vsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-21.5,89.5,9</points>
<connection>
<GID>184</GID>
<name>OUT</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,-21.5,89.5,-21.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-21.5,103.5,10.5</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96,-21.5,103.5,-21.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121,-21.5,121,7.5</points>
<connection>
<GID>192</GID>
<name>OUT</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-21.5,121,-21.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>121 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,-21.5,134,7</points>
<connection>
<GID>194</GID>
<name>OUT</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>125,-21.5,134,-21.5</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>134 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-1.5,73,32.5</points>
<intersection>-1.5 2</intersection>
<intersection>32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,32.5,73,32.5</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,-1.5,75,-1.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-25.5,81,-2.5</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-25.5,125,-25.5</points>
<connection>
<GID>53</GID>
<name>clock_enable</name></connection>
<connection>
<GID>52</GID>
<name>clock_enable</name></connection>
<connection>
<GID>51</GID>
<name>clock_enable</name></connection>
<connection>
<GID>50</GID>
<name>clock_enable</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-153.405,74.6945,177.397,-91.6561</PageViewport>
<gate>
<ID>193</ID>
<type>DE_TO</type>
<position>-15.5,-16</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q3_1</lparam></gate>
<gate>
<ID>195</ID>
<type>DE_TO</type>
<position>-5.5,-16</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q3_0</lparam></gate>
<gate>
<ID>197</ID>
<type>DE_TO</type>
<position>-28,-16</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q3_2</lparam></gate>
<gate>
<ID>199</ID>
<type>DE_TO</type>
<position>-41,-16</position>
<input>
<ID>IN_0</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q3_3</lparam></gate>
<gate>
<ID>200</ID>
<type>AE_OR2</type>
<position>121.5,12</position>
<input>
<ID>IN_0</ID>180 </input>
<input>
<ID>IN_1</ID>179 </input>
<output>
<ID>OUT</ID>191 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_TOGGLE</type>
<position>-46.5,-16</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>202</ID>
<type>AA_TOGGLE</type>
<position>80.5,29.5</position>
<output>
<ID>OUT_0</ID>164 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>203</ID>
<type>AA_TOGGLE</type>
<position>-33,-16</position>
<output>
<ID>OUT_0</ID>150 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>204</ID>
<type>AE_SMALL_INVERTER</type>
<position>57,34.5</position>
<input>
<ID>IN_0</ID>173 </input>
<output>
<ID>OUT_0</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>205</ID>
<type>BE_NOR2</type>
<position>25.5,-86</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>206</ID>
<type>AE_SMALL_INVERTER</type>
<position>78.5,27</position>
<input>
<ID>IN_0</ID>172 </input>
<output>
<ID>OUT_0</ID>165 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_AND2</type>
<position>79.5,21.5</position>
<input>
<ID>IN_0</ID>164 </input>
<input>
<ID>IN_1</ID>165 </input>
<output>
<ID>OUT</ID>178 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_AND2</type>
<position>118,18</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>175 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_TOGGLE</type>
<position>95.5,29</position>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_TOGGLE</type>
<position>110.5,29</position>
<output>
<ID>OUT_0</ID>167 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_TOGGLE</type>
<position>124.5,29.5</position>
<output>
<ID>OUT_0</ID>166 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>212</ID>
<type>AE_SMALL_INVERTER</type>
<position>93.5,27</position>
<input>
<ID>IN_0</ID>172 </input>
<output>
<ID>OUT_0</ID>171 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>213</ID>
<type>AE_SMALL_INVERTER</type>
<position>108.5,27.5</position>
<input>
<ID>IN_0</ID>172 </input>
<output>
<ID>OUT_0</ID>170 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>214</ID>
<type>AE_OR2</type>
<position>91,15.5</position>
<input>
<ID>IN_0</ID>174 </input>
<input>
<ID>IN_1</ID>176 </input>
<output>
<ID>OUT</ID>189 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>AE_SMALL_INVERTER</type>
<position>122,27.5</position>
<input>
<ID>IN_0</ID>172 </input>
<output>
<ID>OUT_0</ID>169 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>216</ID>
<type>DA_FROM</type>
<position>55,44</position>
<input>
<ID>IN_0</ID>173 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID /Load</lparam></gate>
<gate>
<ID>217</ID>
<type>AA_AND2</type>
<position>86.5,21.5</position>
<input>
<ID>IN_0</ID>184 </input>
<input>
<ID>IN_1</ID>175 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_AND2</type>
<position>104,19</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>175 </input>
<output>
<ID>OUT</ID>182 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>219</ID>
<type>AA_AND2</type>
<position>110.5,20</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>170 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_AND2</type>
<position>75.5,37.5</position>
<input>
<ID>IN_0</ID>175 </input>
<input>
<ID>IN_1</ID>173 </input>
<output>
<ID>OUT</ID>172 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND2</type>
<position>94.5,21.5</position>
<input>
<ID>IN_0</ID>168 </input>
<input>
<ID>IN_1</ID>171 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_AND2</type>
<position>123.5,21</position>
<input>
<ID>IN_0</ID>166 </input>
<input>
<ID>IN_1</ID>169 </input>
<output>
<ID>OUT</ID>180 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>223</ID>
<type>AA_AND2</type>
<position>73.5,21</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>175 </input>
<output>
<ID>OUT</ID>177 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>224</ID>
<type>AE_OR2</type>
<position>77,14</position>
<input>
<ID>IN_0</ID>178 </input>
<input>
<ID>IN_1</ID>177 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>225</ID>
<type>AE_OR2</type>
<position>108.5,12.5</position>
<input>
<ID>IN_0</ID>181 </input>
<input>
<ID>IN_1</ID>182 </input>
<output>
<ID>OUT</ID>190 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>AE_OR2</type>
<position>62,11.5</position>
<input>
<ID>IN_0</ID>187 </input>
<input>
<ID>IN_1</ID>186 </input>
<output>
<ID>OUT</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_TOGGLE</type>
<position>-18.5,22</position>
<output>
<ID>OUT_0</ID>192 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>229</ID>
<type>AE_SMALL_INVERTER</type>
<position>-42,27</position>
<input>
<ID>IN_0</ID>197 </input>
<output>
<ID>OUT_0</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>230</ID>
<type>AE_SMALL_INVERTER</type>
<position>-20.5,19.5</position>
<input>
<ID>IN_0</ID>196 </input>
<output>
<ID>OUT_0</ID>193 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>231</ID>
<type>AA_AND2</type>
<position>-19.5,14</position>
<input>
<ID>IN_0</ID>192 </input>
<input>
<ID>IN_1</ID>193 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>232</ID>
<type>AA_TOGGLE</type>
<position>-3.5,21.5</position>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>233</ID>
<type>AE_SMALL_INVERTER</type>
<position>-5.5,19.5</position>
<input>
<ID>IN_0</ID>196 </input>
<output>
<ID>OUT_0</ID>195 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>234</ID>
<type>AE_OR2</type>
<position>-8,8</position>
<input>
<ID>IN_0</ID>198 </input>
<input>
<ID>IN_1</ID>200 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>235</ID>
<type>DA_FROM</type>
<position>-44,36.5</position>
<input>
<ID>IN_0</ID>197 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID /Load</lparam></gate>
<gate>
<ID>236</ID>
<type>AA_AND2</type>
<position>-12.5,14</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>199 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>AA_AND2</type>
<position>-23.5,30</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>197 </input>
<output>
<ID>OUT</ID>196 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>238</ID>
<type>AA_AND2</type>
<position>-4.5,14</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>195 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>239</ID>
<type>AA_AND2</type>
<position>-25.5,13.5</position>
<input>
<ID>IN_0</ID>208 </input>
<input>
<ID>IN_1</ID>199 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>AE_OR2</type>
<position>-22,6.5</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>201 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>241</ID>
<type>AE_OR2</type>
<position>-37,4</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>204 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_LABEL</type>
<position>-18.5,26.5</position>
<gparam>LABEL_TEXT Q3_1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>AA_LABEL</type>
<position>-3,26.5</position>
<gparam>LABEL_TEXT Q3_0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>246</ID>
<type>AA_LABEL</type>
<position>80.5,36</position>
<gparam>LABEL_TEXT Q2_3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>AA_LABEL</type>
<position>92,36</position>
<gparam>LABEL_TEXT Q2_2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>248</ID>
<type>AA_LABEL</type>
<position>108,36.5</position>
<gparam>LABEL_TEXT Q2_1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>249</ID>
<type>AA_LABEL</type>
<position>123.5,36.5</position>
<gparam>LABEL_TEXT Q2_0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>-50,-32</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID H_change</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_AND3</type>
<position>-43.5,-30</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>199 </input>
<input>
<ID>IN_2</ID>50 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>89</ID>
<type>BA_NAND2</type>
<position>-288,-74.5</position>
<input>
<ID>IN_1</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>BE_NOR2</type>
<position>55,-87.5</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>152 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>111</ID>
<type>AE_SMALL_INVERTER</type>
<position>11.5,-79</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>115</ID>
<type>AE_SMALL_INVERTER</type>
<position>47.5,-83.5</position>
<input>
<ID>IN_0</ID>90 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>121</ID>
<type>AF_DFF_LOW</type>
<position>69.5,-23.5</position>
<input>
<ID>IN_0</ID>188 </input>
<output>
<ID>OUTINV_0</ID>107 </output>
<output>
<ID>OUT_0</ID>100 </output>
<input>
<ID>clear</ID>155 </input>
<input>
<ID>clock</ID>118 </input>
<input>
<ID>clock_enable</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>122</ID>
<type>AF_DFF_LOW</type>
<position>84,-23.5</position>
<input>
<ID>IN_0</ID>189 </input>
<output>
<ID>OUTINV_0</ID>106 </output>
<output>
<ID>OUT_0</ID>103 </output>
<input>
<ID>clear</ID>155 </input>
<input>
<ID>clock</ID>118 </input>
<input>
<ID>clock_enable</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>123</ID>
<type>AF_DFF_LOW</type>
<position>98,-23.5</position>
<input>
<ID>IN_0</ID>190 </input>
<output>
<ID>OUTINV_0</ID>101 </output>
<output>
<ID>OUT_0</ID>104 </output>
<input>
<ID>clear</ID>155 </input>
<input>
<ID>clock</ID>118 </input>
<input>
<ID>clock_enable</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>124</ID>
<type>AF_DFF_LOW</type>
<position>113,-23.5</position>
<input>
<ID>IN_0</ID>191 </input>
<output>
<ID>OUTINV_0</ID>102 </output>
<output>
<ID>OUT_0</ID>105 </output>
<input>
<ID>clear</ID>155 </input>
<input>
<ID>clock</ID>118 </input>
<input>
<ID>clock_enable</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_AND3</type>
<position>78.5,-43</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>104 </input>
<input>
<ID>IN_2</ID>103 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_AND3</type>
<position>72,-43</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>101 </input>
<input>
<ID>IN_2</ID>100 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_AND3</type>
<position>89,-43</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>104 </input>
<input>
<ID>IN_2</ID>106 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_AND3</type>
<position>95.5,-43</position>
<input>
<ID>IN_0</ID>101 </input>
<input>
<ID>IN_1</ID>103 </input>
<input>
<ID>IN_2</ID>107 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_AND3</type>
<position>102,-43</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>103 </input>
<input>
<ID>IN_2</ID>107 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_AND3</type>
<position>112.5,-43</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>101 </input>
<input>
<ID>IN_2</ID>107 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>131</ID>
<type>AA_AND2</type>
<position>118,-43</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>114 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>132</ID>
<type>AE_OR2</type>
<position>74,-50</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>133</ID>
<type>AE_OR3</type>
<position>95.5,-50</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>110 </input>
<input>
<ID>IN_2</ID>111 </input>
<output>
<ID>OUT</ID>184 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>134</ID>
<type>AE_OR2</type>
<position>115.5,-49.5</position>
<input>
<ID>IN_0</ID>114 </input>
<input>
<ID>IN_1</ID>113 </input>
<output>
<ID>OUT</ID>183 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>DE_TO</type>
<position>75,-2.5</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q2_3</lparam></gate>
<gate>
<ID>136</ID>
<type>DE_TO</type>
<position>89,-2.5</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q2_2</lparam></gate>
<gate>
<ID>137</ID>
<type>DE_TO</type>
<position>102.5,-3</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q2_1</lparam></gate>
<gate>
<ID>138</ID>
<type>DE_TO</type>
<position>116.5,-3</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q2_0</lparam></gate>
<gate>
<ID>139</ID>
<type>AA_AND2</type>
<position>-316,-65.5</position>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_AND2</type>
<position>-291,-72.5</position>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>141</ID>
<type>AA_AND2</type>
<position>-300,-39.5</position>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_AND2</type>
<position>-292,-79</position>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>DA_FROM</type>
<position>40.5,-83</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /MR2</lparam></gate>
<gate>
<ID>148</ID>
<type>DA_FROM</type>
<position>57,-11</position>
<input>
<ID>IN_0</ID>118 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_AND2</type>
<position>54.5,-26</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>175 </input>
<output>
<ID>OUT</ID>186 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>154</ID>
<type>DA_FROM</type>
<position>-32,-21</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Clk</lparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>45.5,-27</position>
<input>
<ID>IN_0</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>160</ID>
<type>AE_SMALL_INVERTER</type>
<position>-272,-62</position>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>162</ID>
<type>AA_TOGGLE</type>
<position>-80,-8.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>164</ID>
<type>AF_DFF_LOW</type>
<position>-24,-31.5</position>
<input>
<ID>IN_0</ID>205 </input>
<output>
<ID>OUTINV_0</ID>129 </output>
<output>
<ID>OUT_0</ID>153 </output>
<input>
<ID>clear</ID>154 </input>
<input>
<ID>clock</ID>145 </input>
<input>
<ID>clock_enable</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>166</ID>
<type>AF_DFF_LOW</type>
<position>-8,-31.5</position>
<input>
<ID>IN_0</ID>206 </input>
<output>
<ID>OUTINV_0</ID>131 </output>
<output>
<ID>OUT_0</ID>130 </output>
<input>
<ID>clear</ID>154 </input>
<input>
<ID>clock</ID>145 </input>
<input>
<ID>clock_enable</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>168</ID>
<type>AA_AND2</type>
<position>-20,-46.5</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>208 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_AND2</type>
<position>-3,-46.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_AND2</type>
<position>-315.5,-40.5</position>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_AND2</type>
<position>-292.5,-57.5</position>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>DA_FROM</type>
<position>2,-78.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /MR3</lparam></gate>
<gate>
<ID>178</ID>
<type>AE_SMALL_INVERTER</type>
<position>-308,-52</position>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>180</ID>
<type>AA_AND2</type>
<position>29.5,-72.5</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>153 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>181</ID>
<type>DA_FROM</type>
<position>46,-25</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID H_change</lparam></gate>
<gate>
<ID>183</ID>
<type>AA_AND2</type>
<position>-315.5,-59.5</position>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_AND2</type>
<position>-301.5,-66.5</position>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_AND2</type>
<position>0,-6</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>DA_FROM</type>
<position>-52,-30</position>
<input>
<ID>IN_0</ID>199 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID CE</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_AND2</type>
<position>-285,-44</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>-20.5,17,-20.5,17.5</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,17,-3.5,19.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,17,-5.5,17.5</points>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>-23.5,24,-23.5,27</points>
<connection>
<GID>237</GID>
<name>OUT</name></connection>
<intersection>24 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-23.5,24,-5.5,24</points>
<intersection>-23.5 1</intersection>
<intersection>-20.5 10</intersection>
<intersection>-5.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-5.5,21.5,-5.5,24</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>24 2</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>-20.5,21.5,-20.5,24</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>24 2</intersection></vsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,34,-24.5,34</points>
<intersection>-27.5 5</intersection>
<intersection>-24.5 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-27.5,34,-27.5,36.5</points>
<intersection>34 1</intersection>
<intersection>36.5 8</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>-24.5,33,-24.5,34</points>
<connection>
<GID>237</GID>
<name>IN_1</name></connection>
<intersection>34 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-44,36.5,-27.5,36.5</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>-44 9</intersection>
<intersection>-27.5 5</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-44,27,-44,36.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>36.5 8</intersection></vsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7,11,-4.5,11</points>
<connection>
<GID>238</GID>
<name>OUT</name></connection>
<connection>
<GID>234</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>-35,26.5,-35,33</points>
<intersection>26.5 4</intersection>
<intersection>28.5 10</intersection>
<intersection>33 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-35,33,-22.5,33</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>-35 2</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-35,26.5,-13.5,26.5</points>
<intersection>-35 2</intersection>
<intersection>-26.5 9</intersection>
<intersection>-13.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-13.5,17,-13.5,26.5</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<intersection>26.5 4</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-26.5,16.5,-26.5,26.5</points>
<connection>
<GID>239</GID>
<name>IN_1</name></connection>
<intersection>26.5 4</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-46.5,28.5,-35,28.5</points>
<intersection>-46.5 20</intersection>
<intersection>-35 2</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>-50,-29.5,-46.5,-29.5</points>
<intersection>-50 21</intersection>
<intersection>-46.5 20</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>-46.5,-30,-46.5,28.5</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>-29.5 12</intersection>
<intersection>28.5 10</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>-50,-30,-50,-29.5</points>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>-29.5 12</intersection></vsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12.5,11,-9,11</points>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<connection>
<GID>234</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23,9.5,-23,10</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<intersection>10 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-25.5,10,-25.5,10.5</points>
<connection>
<GID>239</GID>
<name>OUT</name></connection>
<intersection>10 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-25.5,10,-23,10</points>
<intersection>-25.5 1</intersection>
<intersection>-23 0</intersection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,10,-19.5,11</points>
<connection>
<GID>231</GID>
<name>OUT</name></connection>
<intersection>10 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-21,9.5,-21,10</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>10 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-21,10,-19.5,10</points>
<intersection>-21 1</intersection>
<intersection>-19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,5,-40,27</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40,-30,-40,3</points>
<connection>
<GID>241</GID>
<name>IN_1</name></connection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-40.5,-30,-40,-30</points>
<connection>
<GID>81</GID>
<name>OUT</name></connection>
<intersection>-40 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-29.5,-22,3.5</points>
<connection>
<GID>240</GID>
<name>OUT</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27,-29.5,-22,-29.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,-29.5,-8,5</points>
<connection>
<GID>234</GID>
<name>OUT</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11,-29.5,-8,-29.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>-8 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,-16,-11.5,17</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>-16 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-3,-49.5,-3,-16</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-11.5,-16,-3,-16</points>
<intersection>-11.5 0</intersection>
<intersection>-3 1</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24.5,-16.5,-24.5,16.5</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>-16.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-20,-49.5,-20,-16.5</points>
<connection>
<GID>168</GID>
<name>OUT</name></connection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-24.5,-16.5,-20,-16.5</points>
<intersection>-24.5 0</intersection>
<intersection>-20 1</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-48,-32,-46.5,-32</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<connection>
<GID>81</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54,-28,-54,-6</points>
<intersection>-28 1</intersection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-54,-28,-46.5,-28</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>-54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-54,-6,-3,-6</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<intersection>-54 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-291,-75.5,-291,-75.5</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<connection>
<GID>140</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-44.5,-16,-43,-16</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-79,6.5,-78.5</points>
<intersection>-79 1</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-79,9.5,-79</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,-78.5,6.5,-78.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-83,24.5,-79</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-79,24.5,-79</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44,-83.5,44,-83</points>
<intersection>-83.5 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,-83.5,45.5,-83.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42.5,-83,44,-83</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>44 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-86.5,50.5,-83.5</points>
<intersection>-86.5 1</intersection>
<intersection>-83.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-86.5,52,-86.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-83.5,50.5,-83.5</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-29.5,73.5,-21.5</points>
<intersection>-29.5 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-21.5,73.5,-21.5</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<intersection>72.5 4</intersection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-29.5,73.5,-29.5</points>
<intersection>70 3</intersection>
<intersection>73.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70,-40,70,-29.5</points>
<connection>
<GID>126</GID>
<name>IN_2</name></connection>
<intersection>-29.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>72.5,-21.5,72.5,-2.5</points>
<intersection>-21.5 1</intersection>
<intersection>-5 6</intersection>
<intersection>-2.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>72.5,-2.5,73,-2.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>72.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>3,-5,72.5,-5</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>72.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-40,72,-37.5</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-37.5,112.5,-37.5</points>
<intersection>72 0</intersection>
<intersection>97.5 3</intersection>
<intersection>101 2</intersection>
<intersection>112.5 4</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>101,-37.5,101,-24.5</points>
<connection>
<GID>123</GID>
<name>OUTINV_0</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>97.5,-40,97.5,-37.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>112.5,-40,112.5,-37.5</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>-37.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74,-39,127.5,-39</points>
<intersection>74 26</intersection>
<intersection>104 3</intersection>
<intersection>119 4</intersection>
<intersection>127.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>127.5,-39,127.5,-10.5</points>
<intersection>-39 1</intersection>
<intersection>-24.5 31</intersection>
<intersection>-10.5 29</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>104,-40,104,-39</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>119,-40,119,-39</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment>
<vsegment>
<ID>26</ID>
<points>74,-40,74,-39</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>119,-10.5,127.5,-10.5</points>
<intersection>119 32</intersection>
<intersection>127.5 2</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>116,-24.5,127.5,-24.5</points>
<connection>
<GID>124</GID>
<name>OUTINV_0</name></connection>
<intersection>127.5 2</intersection></hsegment>
<vsegment>
<ID>32</ID>
<points>119,-10.5,119,21</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>-10.5 29</intersection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-31,88,-21.5</points>
<intersection>-31 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-21.5,88,-21.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>87 9</intersection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76.5,-31,102,-31</points>
<intersection>76.5 3</intersection>
<intersection>88 0</intersection>
<intersection>95.5 6</intersection>
<intersection>102 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>76.5,-69.5,76.5,-31</points>
<connection>
<GID>125</GID>
<name>IN_2</name></connection>
<intersection>-69.5 10</intersection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>95.5,-40,95.5,-31</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>102,-40,102,-31</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>-31 2</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>87,-21.5,87,-2.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>30.5,-69.5,76.5,-69.5</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>76.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-32,102.5,-21.5</points>
<intersection>-32 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-21.5,102.5,-21.5</points>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<intersection>100.5 7</intersection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78.5,-32,117,-32</points>
<intersection>78.5 3</intersection>
<intersection>89 4</intersection>
<intersection>102.5 0</intersection>
<intersection>117 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>78.5,-40,78.5,-32</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>89,-40,89,-32</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>117,-40,117,-32</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>-32 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>100.5,-21.5,100.5,-3</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>-21.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-33,118,-21.5</points>
<intersection>-33 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>114.5,-21.5,118,-21.5</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>114.5 6</intersection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3,-33,118,-33</points>
<intersection>3 8</intersection>
<intersection>80.5 3</intersection>
<intersection>91 4</intersection>
<intersection>114.5 5</intersection>
<intersection>118 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>80.5,-40,80.5,-33</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>-33 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>91,-40,91,-33</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>-33 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>114.5,-40,114.5,-33</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-33 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>114.5,-21.5,114.5,-3</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>3,-33,3,-7</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>-33 2</intersection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-40,87,-24.5</points>
<connection>
<GID>122</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>127</GID>
<name>IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,-40,93.5,-35.5</points>
<connection>
<GID>128</GID>
<name>IN_2</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-35.5,110.5,-35.5</points>
<intersection>72.5 2</intersection>
<intersection>93.5 0</intersection>
<intersection>100 4</intersection>
<intersection>110.5 6</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>72.5,-35.5,72.5,-24.5</points>
<connection>
<GID>121</GID>
<name>OUTINV_0</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>100,-40,100,-35.5</points>
<connection>
<GID>129</GID>
<name>IN_2</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>110.5,-40,110.5,-35.5</points>
<connection>
<GID>130</GID>
<name>IN_2</name></connection>
<intersection>-35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-47,75,-46.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>78.5,-46.5,78.5,-46</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>75,-46.5,78.5,-46.5</points>
<intersection>75 0</intersection>
<intersection>78.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-47,73,-46.5</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>72,-46.5,72,-46</points>
<connection>
<GID>126</GID>
<name>OUT</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>72,-46.5,73,-46.5</points>
<intersection>72 1</intersection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-47,95.5,-46</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<connection>
<GID>128</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-46.5,89,-46</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>93.5,-47,93.5,-46.5</points>
<connection>
<GID>133</GID>
<name>IN_2</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>89,-46.5,93.5,-46.5</points>
<intersection>89 0</intersection>
<intersection>93.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-46.5,102,-46</points>
<connection>
<GID>129</GID>
<name>OUT</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>97.5,-47,97.5,-46.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-46.5,102,-46.5</points>
<intersection>97.5 1</intersection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-46.5,114.5,-46</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>112.5,-46,114.5,-46</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-46.5,116.5,-46</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>-46 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-46,118,-46</points>
<connection>
<GID>131</GID>
<name>OUT</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>59,-11,108.5,-11</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>65.5 9</intersection>
<intersection>80 8</intersection>
<intersection>94 7</intersection>
<intersection>108.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>108.5,-23.5,108.5,-11</points>
<intersection>-23.5 17</intersection>
<intersection>-11 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>94,-23.5,94,-11</points>
<intersection>-23.5 12</intersection>
<intersection>-11 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>80,-23.5,80,-11</points>
<intersection>-23.5 11</intersection>
<intersection>-11 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>65.5,-23.5,65.5,-11</points>
<intersection>-23.5 16</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>80,-23.5,81,-23.5</points>
<connection>
<GID>122</GID>
<name>clock</name></connection>
<intersection>80 8</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>94,-23.5,95,-23.5</points>
<connection>
<GID>123</GID>
<name>clock</name></connection>
<intersection>94 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>65.5,-23.5,66.5,-23.5</points>
<connection>
<GID>121</GID>
<name>clock</name></connection>
<intersection>65.5 9</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>108.5,-23.5,110,-23.5</points>
<connection>
<GID>124</GID>
<name>clock</name></connection>
<intersection>108.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>65.5,-29,110,-29</points>
<intersection>65.5 8</intersection>
<intersection>81 7</intersection>
<intersection>95 10</intersection>
<intersection>110 12</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>81,-29,81,-25.5</points>
<connection>
<GID>122</GID>
<name>clock_enable</name></connection>
<intersection>-29 5</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>65.5,-29,65.5,11.5</points>
<intersection>-29 5</intersection>
<intersection>-25.5 15</intersection>
<intersection>11.5 16</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>95,-29,95,-25.5</points>
<connection>
<GID>123</GID>
<name>clock_enable</name></connection>
<intersection>-29 5</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>110,-29,110,-25.5</points>
<connection>
<GID>124</GID>
<name>clock_enable</name></connection>
<intersection>-29 5</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>65.5,-25.5,66.5,-25.5</points>
<connection>
<GID>121</GID>
<name>clock_enable</name></connection>
<intersection>65.5 8</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>65,11.5,65.5,11.5</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<intersection>65.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-43.5,-21,-32.5</points>
<connection>
<GID>164</GID>
<name>OUTINV_0</name></connection>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>-43.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-21,-43.5,-4,-43.5</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-41,-4,-29.5</points>
<intersection>-41 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-29.5,-4,-29.5</points>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<intersection>-5 5</intersection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19,-41,-4,-41</points>
<intersection>-19 3</intersection>
<intersection>-4 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-19,-43.5,-19,-41</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>-41 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-5,-29.5,-5,-21</points>
<intersection>-29.5 1</intersection>
<intersection>-21 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-7.5,-21,-5,-21</points>
<intersection>-7.5 7</intersection>
<intersection>-5 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-7.5,-21,-7.5,-16</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>-21 6</intersection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-43.5,-2,-32.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5,-32.5,-2,-32.5</points>
<connection>
<GID>166</GID>
<name>OUTINV_0</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-25,51.5,-25</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<connection>
<GID>181</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30,-21,-12.5,-21</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>-28 5</intersection>
<intersection>-12.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-12.5,-31.5,-12.5,-21</points>
<intersection>-31.5 6</intersection>
<intersection>-21 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-28,-31.5,-28,-21</points>
<intersection>-31.5 7</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-12.5,-31.5,-11,-31.5</points>
<connection>
<GID>166</GID>
<name>clock</name></connection>
<intersection>-12.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-28,-31.5,-27,-31.5</points>
<connection>
<GID>164</GID>
<name>clock</name></connection>
<intersection>-28 5</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-32,-38.5,-11,-38.5</points>
<intersection>-32 5</intersection>
<intersection>-11 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-11,-38.5,-11,-33.5</points>
<connection>
<GID>166</GID>
<name>clock_enable</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-32,-38.5,-32,4</points>
<intersection>-38.5 1</intersection>
<intersection>-33.5 10</intersection>
<intersection>4 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-34,4,-32,4</points>
<connection>
<GID>241</GID>
<name>OUT</name></connection>
<intersection>-32 5</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-32,-33.5,-27,-33.5</points>
<connection>
<GID>164</GID>
<name>clock_enable</name></connection>
<intersection>-32 5</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-31,-16,-30,-16</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-88.5,29.5,-75.5</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<intersection>-88.5 4</intersection>
<intersection>-79 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>26.5,-83,26.5,-79</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>-79 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-79,29.5,-79</points>
<intersection>26.5 1</intersection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>29.5,-88.5,52,-88.5</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,-69.5,-20.5,-16</points>
<intersection>-69.5 4</intersection>
<intersection>-29.5 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-29.5,-20.5,-29.5</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>-20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-20.5,-16,-17.5,-16</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>-20.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-20.5,-69.5,28.5,-69.5</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>-20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-91,-42.5,-35.5</points>
<intersection>-91 2</intersection>
<intersection>-35.5 3</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>25.5,-91,25.5,-89</points>
<connection>
<GID>205</GID>
<name>OUT</name></connection>
<intersection>-91 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-42.5,-91,25.5,-91</points>
<intersection>-42.5 0</intersection>
<intersection>25.5 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-42.5,-35.5,-8,-35.5</points>
<connection>
<GID>166</GID>
<name>clear</name></connection>
<connection>
<GID>164</GID>
<name>clear</name></connection>
<intersection>-42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<hsegment>
<ID>4</ID>
<points>58,-27.5,113,-27.5</points>
<connection>
<GID>121</GID>
<name>clear</name></connection>
<connection>
<GID>124</GID>
<name>clear</name></connection>
<connection>
<GID>123</GID>
<name>clear</name></connection>
<connection>
<GID>122</GID>
<name>clear</name></connection>
<intersection>58 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>58,-87.5,58,-27.5</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>-27.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,24.5,80.5,27.5</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>4</ID>
<points>78.5,24.5,78.5,25</points>
<connection>
<GID>207</GID>
<name>IN_1</name></connection>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,24,124.5,27.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<connection>
<GID>211</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,23,111.5,27</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>27 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>110.5,27,111.5,27</points>
<connection>
<GID>210</GID>
<name>OUT_0</name></connection>
<intersection>111.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,24.5,95.5,27</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,24,122.5,24.5</points>
<connection>
<GID>222</GID>
<name>IN_1</name></connection>
<intersection>24.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>122,24.5,122,25.5</points>
<connection>
<GID>215</GID>
<name>OUT_0</name></connection>
<intersection>24.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>122,24.5,122.5,24.5</points>
<intersection>122 1</intersection>
<intersection>122.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>6</ID>
<points>109.5,23,109.5,25.5</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>25.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>108.5,25.5,109.5,25.5</points>
<connection>
<GID>213</GID>
<name>OUT_0</name></connection>
<intersection>109.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,24.5,93.5,25</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>1</ID>
<points>75.5,31.5,75.5,34.5</points>
<connection>
<GID>220</GID>
<name>OUT</name></connection>
<intersection>31.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>75.5,31.5,122,31.5</points>
<intersection>75.5 1</intersection>
<intersection>78.5 10</intersection>
<intersection>93.5 4</intersection>
<intersection>108.5 6</intersection>
<intersection>122 8</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>93.5,29,93.5,31.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>31.5 2</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>108.5,29.5,108.5,31.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>31.5 2</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>122,29.5,122,31.5</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>31.5 2</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>78.5,29,78.5,31.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>31.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71.5,41.5,74.5,41.5</points>
<intersection>71.5 5</intersection>
<intersection>74.5 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>71.5,41.5,71.5,44</points>
<intersection>41.5 1</intersection>
<intersection>44 8</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>74.5,40.5,74.5,41.5</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<intersection>41.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>55,44,71.5,44</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>55 9</intersection>
<intersection>71.5 5</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>55,34.5,55,44</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>44 8</intersection></vsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>92,18.5,94.5,18.5</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<connection>
<GID>214</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>2</ID>
<points>64,34,64,40.5</points>
<intersection>34 4</intersection>
<intersection>36.5 10</intersection>
<intersection>40.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>64,40.5,76.5,40.5</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>64 2</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>64,34,117,34</points>
<intersection>64 2</intersection>
<intersection>72.5 9</intersection>
<intersection>85.5 5</intersection>
<intersection>103 8</intersection>
<intersection>117 7</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>85.5,24.5,85.5,34</points>
<connection>
<GID>217</GID>
<name>IN_1</name></connection>
<intersection>34 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>117,21,117,34</points>
<connection>
<GID>208</GID>
<name>IN_1</name></connection>
<intersection>34 4</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>103,22,103,34</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<intersection>34 4</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>72.5,24,72.5,34</points>
<connection>
<GID>223</GID>
<name>IN_1</name></connection>
<intersection>34 4</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>51.5,36.5,64,36.5</points>
<intersection>51.5 13</intersection>
<intersection>64 2</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>47.5,-27.5,51.5,-27.5</points>
<intersection>47.5 14</intersection>
<intersection>51.5 13</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>51.5,-27.5,51.5,36.5</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>-27.5 12</intersection>
<intersection>36.5 10</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>47.5,-27.5,47.5,-27</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>-27.5 12</intersection></vsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,18.5,90,18.5</points>
<connection>
<GID>217</GID>
<name>OUT</name></connection>
<connection>
<GID>214</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,17,76,17.5</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<intersection>17.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>73.5,17.5,73.5,18</points>
<connection>
<GID>223</GID>
<name>OUT</name></connection>
<intersection>17.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>73.5,17.5,76,17.5</points>
<intersection>73.5 1</intersection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,17.5,79.5,18.5</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<intersection>17.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>78,17,78,17.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>17.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>78,17.5,79.5,17.5</points>
<intersection>78 1</intersection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118,15,120.5,15</points>
<connection>
<GID>208</GID>
<name>OUT</name></connection>
<connection>
<GID>200</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,16.5,123.5,18</points>
<connection>
<GID>222</GID>
<name>OUT</name></connection>
<intersection>16.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>122.5,15,122.5,16.5</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>16.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>122.5,16.5,123.5,16.5</points>
<intersection>122.5 1</intersection>
<intersection>123.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,16,110.5,17</points>
<connection>
<GID>219</GID>
<name>OUT</name></connection>
<intersection>16 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>109.5,15.5,109.5,16</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>109.5,16,110.5,16</points>
<intersection>109.5 1</intersection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,15.5,104,16</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<intersection>15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>104,15.5,107.5,15.5</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-52.5,115.5,-15</points>
<connection>
<GID>134</GID>
<name>OUT</name></connection>
<intersection>-15 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>105,-15,105,22</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>105,-15,115.5,-15</points>
<intersection>105 1</intersection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-53,95.5,-14</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<intersection>-14 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>87.5,-14,87.5,24.5</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-14,95.5,-14</points>
<intersection>87.5 1</intersection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-14.5,74.5,24</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>74,-53,74,-14.5</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>74,-14.5,74.5,-14.5</points>
<intersection>74 1</intersection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-26,58.5,10.5</points>
<intersection>-26 2</intersection>
<intersection>10.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-26,58.5,-26</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>58.5,10.5,59,10.5</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,12.5,59,34.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-21.5,77,11</points>
<connection>
<GID>224</GID>
<name>OUT</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-21.5,77,-21.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>77 0</intersection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-21.5,91,12.5</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-21.5,91,-21.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>91 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108.5,-21.5,108.5,9.5</points>
<connection>
<GID>225</GID>
<name>OUT</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95,-21.5,108.5,-21.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>108.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-21.5,121.5,9</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>110,-21.5,121.5,-21.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>121.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18.5,17,-18.5,20</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<connection>
<GID>228</GID>
<name>OUT_0</name></connection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,1660.22,1394,959.221</PageViewport></page 3>
<page 4>
<PageViewport>0,1660.22,1394,959.221</PageViewport></page 4>
<page 5>
<PageViewport>0,1660.22,1394,959.221</PageViewport></page 5>
<page 6>
<PageViewport>0,1660.22,1394,959.221</PageViewport></page 6>
<page 7>
<PageViewport>0,1660.22,1394,959.221</PageViewport></page 7>
<page 8>
<PageViewport>0,1660.22,1394,959.221</PageViewport></page 8>
<page 9>
<PageViewport>0,1660.22,1394,959.221</PageViewport></page 9></circuit>