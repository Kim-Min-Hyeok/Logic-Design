<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-81.36,69.7332,506.07,-225.668</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>9.5,-15.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>9.5,-18</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>9.5,-20.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>9.5,-23</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>5</ID>
<type>AI_XOR3</type>
<position>19.5,-25.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>6</ID>
<type>AI_XOR3</type>
<position>19.5,-32</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>7</ID>
<type>AI_XOR3</type>
<position>19.5,-38.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>7 </input>
<input>
<ID>IN_2</ID>6 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>28.5,-15.5</position>
<input>
<ID>N_in0</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>GA_LED</type>
<position>28.5,-18</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>28.5,-20.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>GA_LED</type>
<position>28.5,-25.5</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>28.5,-32</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>28.5,-38.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>6,-15</position>
<gparam>LABEL_TEXT m1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>6,-17.5</position>
<gparam>LABEL_TEXT m2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>6,-20</position>
<gparam>LABEL_TEXT m3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>6,-22.5</position>
<gparam>LABEL_TEXT m4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>GA_LED</type>
<position>28.5,-23</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>31.5,-24.5</position>
<gparam>LABEL_TEXT p1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>31.5,-31</position>
<gparam>LABEL_TEXT p2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>31.5,-37.5</position>
<gparam>LABEL_TEXT p3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>19.5,-8.5</position>
<gparam>LABEL_TEXT Encoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AI_XOR2</type>
<position>106,-13</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AI_XOR2</type>
<position>106,-17.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>AI_XOR2</type>
<position>106,-22</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>AI_XOR2</type>
<position>106,-26.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>AI_XOR2</type>
<position>106,-31</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>AI_XOR2</type>
<position>106,-35.5</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AI_XOR2</type>
<position>106,-40</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>GA_LED</type>
<position>114,-13</position>
<input>
<ID>N_in0</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>114,-17.5</position>
<input>
<ID>N_in0</ID>71 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>114,-22</position>
<input>
<ID>N_in0</ID>72 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>GA_LED</type>
<position>114,-26.5</position>
<input>
<ID>N_in0</ID>73 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>GA_LED</type>
<position>114,-31</position>
<input>
<ID>N_in0</ID>74 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>GA_LED</type>
<position>114,-35.5</position>
<input>
<ID>N_in0</ID>75 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>114,-40</position>
<input>
<ID>N_in0</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AI_XOR4</type>
<position>68,-17</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>57 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>77 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>88</ID>
<type>AI_XOR4</type>
<position>68,-27</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>59 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>78 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>89</ID>
<type>AI_XOR4</type>
<position>68,-36.5</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>59 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>79 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>90</ID>
<type>BE_DECODER_3x8</type>
<position>89.5,-26</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>61 </input>
<input>
<ID>IN_2</ID>60 </input>
<output>
<ID>OUT_1</ID>63 </output>
<output>
<ID>OUT_2</ID>64 </output>
<output>
<ID>OUT_3</ID>65 </output>
<output>
<ID>OUT_4</ID>66 </output>
<output>
<ID>OUT_5</ID>67 </output>
<output>
<ID>OUT_6</ID>68 </output>
<output>
<ID>OUT_7</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_TOGGLE</type>
<position>38,-15</position>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_TOGGLE</type>
<position>38,-17.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>93</ID>
<type>AA_TOGGLE</type>
<position>38,-20</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>38,-22.5</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_TOGGLE</type>
<position>38,-25</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_TOGGLE</type>
<position>38,-27.5</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_TOGGLE</type>
<position>38,-30</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>75.5,-7</position>
<gparam>LABEL_TEXT Decoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>44,-54.5</position>
<gparam>LABEL_TEXT The pull model is on Page2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-15.5,27.5,-15.5</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>16 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>16,-30,16,-15.5</points>
<intersection>-30 6</intersection>
<intersection>-23.5 7</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>16,-30,16.5,-30</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>16 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>16,-23.5,16.5,-23.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>16 4</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-18,27.5,-18</points>
<connection>
<GID>9</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>14.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14.5,-25.5,14.5,-18</points>
<intersection>-25.5 4</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>14.5,-25.5,16.5,-25.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>14.5 3</intersection>
<intersection>16 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>16,-36.5,16,-25.5</points>
<intersection>-36.5 6</intersection>
<intersection>-25.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>16,-36.5,16.5,-36.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>16 5</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-38.5,27.5,-38.5</points>
<connection>
<GID>13</GID>
<name>N_in0</name></connection>
<connection>
<GID>7</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-32,27.5,-32</points>
<connection>
<GID>12</GID>
<name>N_in0</name></connection>
<connection>
<GID>6</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-25.5,27.5,-25.5</points>
<connection>
<GID>11</GID>
<name>N_in0</name></connection>
<connection>
<GID>5</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-40.5,12,-23</points>
<intersection>-40.5 6</intersection>
<intersection>-34 4</intersection>
<intersection>-27.5 9</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-23,27.5,-23</points>
<connection>
<GID>18</GID>
<name>N_in0</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>12,-34,16.5,-34</points>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>12,-40.5,16.5,-40.5</points>
<connection>
<GID>7</GID>
<name>IN_2</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>12,-27.5,16.5,-27.5</points>
<connection>
<GID>5</GID>
<name>IN_2</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-38.5,13.5,-20.5</points>
<intersection>-38.5 4</intersection>
<intersection>-32 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11.5,-20.5,27.5,-20.5</points>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-32,16.5,-32</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>13.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>13.5,-38.5,16.5,-38.5</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-15,65,-15</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<intersection>50 4</intersection>
<intersection>65 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>50,-24,50,-12</points>
<intersection>-24 5</intersection>
<intersection>-15 1</intersection>
<intersection>-12 10</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>50,-24,65,-24</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>50 4</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>50,-12,103,-12</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>50 4</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>65,-15,65,-14</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>-15 1</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-33.5,52.5,-16</points>
<intersection>-33.5 4</intersection>
<intersection>-17.5 6</intersection>
<intersection>-16.5 10</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-16,65,-16</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52.5,-33.5,65,-33.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>40,-17.5,52.5,-17.5</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>52.5,-16.5,103,-16.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-37.5,56,-18</points>
<intersection>-37.5 5</intersection>
<intersection>-28 3</intersection>
<intersection>-25.5 10</intersection>
<intersection>-22.5 6</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-18,65,-18</points>
<connection>
<GID>87</GID>
<name>IN_2</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>56,-28,65,-28</points>
<connection>
<GID>88</GID>
<name>IN_2</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>56,-37.5,65,-37.5</points>
<connection>
<GID>89</GID>
<name>IN_2</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>40,-22.5,56,-22.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>56,-25.5,103,-25.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-35.5,45.5,-20</points>
<intersection>-35.5 4</intersection>
<intersection>-26 2</intersection>
<intersection>-21 9</intersection>
<intersection>-20 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-26,65,-26</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>45.5,-35.5,65,-35.5</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>40,-20,45.5,-20</points>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>45.5,-21,103,-21</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-27.5,80,-17</points>
<intersection>-27.5 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-27.5,86.5,-27.5</points>
<connection>
<GID>90</GID>
<name>IN_2</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-17,80,-17</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-28.5,79,-27</points>
<intersection>-28.5 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-28.5,86.5,-28.5</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-27,79,-27</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79,-36.5,79,-29.5</points>
<intersection>-36.5 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-29.5,86.5,-29.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>79 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>72,-36.5,79,-36.5</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<intersection>79 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94,-41,94,-28.5</points>
<intersection>-41 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94,-41,103,-41</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>94 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-28.5,94,-28.5</points>
<connection>
<GID>90</GID>
<name>OUT_1</name></connection>
<intersection>94 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-36.5,95,-27.5</points>
<intersection>-36.5 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92.5,-27.5,95,-27.5</points>
<connection>
<GID>90</GID>
<name>OUT_2</name></connection>
<intersection>95 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95,-36.5,103,-36.5</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>95 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-26.5,96.5,-23</points>
<intersection>-26.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96.5,-23,103,-23</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-26.5,96.5,-26.5</points>
<connection>
<GID>90</GID>
<name>OUT_3</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-32,98,-25.5</points>
<intersection>-32 1</intersection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98,-32,103,-32</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>98 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-25.5,98,-25.5</points>
<connection>
<GID>90</GID>
<name>OUT_4</name></connection>
<intersection>98 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-24.5,99.5,-18.5</points>
<intersection>-24.5 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-18.5,103,-18.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-24.5,99.5,-24.5</points>
<connection>
<GID>90</GID>
<name>OUT_5</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-23.5,100.5,-14</points>
<intersection>-23.5 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-14,103,-14</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-23.5,100.5,-23.5</points>
<connection>
<GID>90</GID>
<name>OUT_6</name></connection>
<intersection>100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101.5,-27.5,101.5,-22.5</points>
<intersection>-27.5 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>101.5,-27.5,103,-27.5</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>101.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-22.5,101.5,-22.5</points>
<connection>
<GID>90</GID>
<name>OUT_7</name></connection>
<intersection>101.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-13,113,-13</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<connection>
<GID>80</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-17.5,113,-17.5</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<connection>
<GID>81</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-22,113,-22</points>
<connection>
<GID>75</GID>
<name>OUT</name></connection>
<connection>
<GID>82</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-26.5,113,-26.5</points>
<connection>
<GID>76</GID>
<name>OUT</name></connection>
<connection>
<GID>83</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-31,113,-31</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<connection>
<GID>84</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-35.5,113,-35.5</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<connection>
<GID>85</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-40,113,-40</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<connection>
<GID>86</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-30,48,-25</points>
<intersection>-30 6</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-25,65,-25</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>48 0</intersection>
<intersection>65 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>65,-25,65,-20</points>
<connection>
<GID>87</GID>
<name>IN_3</name></connection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>48,-30,103,-30</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-34.5,43.5,-27.5</points>
<intersection>-34.5 6</intersection>
<intersection>-30 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-30,65,-30</points>
<connection>
<GID>88</GID>
<name>IN_3</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-27.5,43.5,-27.5</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>43.5,-34.5,103,-34.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-39.5,41.5,-30</points>
<intersection>-39.5 1</intersection>
<intersection>-39 6</intersection>
<intersection>-30 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-39.5,65,-39.5</points>
<connection>
<GID>89</GID>
<name>IN_3</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-30,41.5,-30</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>41.5,-39,103,-39</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-79.5777,18.8305,106.289,-74.6362</PageViewport>
<gate>
<ID>100</ID>
<type>AI_XOR2</type>
<position>42.5,-1.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>101</ID>
<type>AI_XOR2</type>
<position>42.5,-6</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AI_XOR2</type>
<position>42.5,-10.5</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>AI_XOR2</type>
<position>42.5,-15</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AI_XOR2</type>
<position>42.5,-19.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>107 </input>
<output>
<ID>OUT</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>105</ID>
<type>AI_XOR2</type>
<position>42.5,-24</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>105 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AI_XOR2</type>
<position>42.5,-28.5</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_TOGGLE</type>
<position>-51,-2.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_TOGGLE</type>
<position>-51,-5</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_TOGGLE</type>
<position>-51,-7.5</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_TOGGLE</type>
<position>-51,-10</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>111</ID>
<type>AI_XOR3</type>
<position>-40.5,-19.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>81 </input>
<input>
<ID>IN_2</ID>82 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>112</ID>
<type>AI_XOR3</type>
<position>-40.5,-26</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>82 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>113</ID>
<type>AI_XOR3</type>
<position>-40.5,-32.5</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>82 </input>
<output>
<ID>OUT</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>-54.5,-2</position>
<gparam>LABEL_TEXT m1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>-54.5,-4.5</position>
<gparam>LABEL_TEXT m2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>-54.5,-7</position>
<gparam>LABEL_TEXT m3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>-54.5,-9.5</position>
<gparam>LABEL_TEXT m4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_TOGGLE</type>
<position>-43,4</position>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_TOGGLE</type>
<position>-40.5,4</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_TOGGLE</type>
<position>-38,4</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_TOGGLE</type>
<position>-35.5,4</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_TOGGLE</type>
<position>-33,4</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_TOGGLE</type>
<position>-30.5,4</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_TOGGLE</type>
<position>-28,4</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>125</ID>
<type>AI_XOR2</type>
<position>-18,-2.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>84 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AI_XOR2</type>
<position>-18,-7</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>85 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>AI_XOR2</type>
<position>-18,-11.5</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>128</ID>
<type>AI_XOR2</type>
<position>-18,-16</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>129</ID>
<type>AI_XOR2</type>
<position>-18,-20.5</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>130</ID>
<type>AI_XOR2</type>
<position>-18,-25</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>131</ID>
<type>AI_XOR2</type>
<position>-18,-29.5</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>132</ID>
<type>AI_XOR4</type>
<position>4.5,-5.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<input>
<ID>IN_2</ID>96 </input>
<input>
<ID>IN_3</ID>97 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>133</ID>
<type>AI_XOR4</type>
<position>4.5,-15.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>98 </input>
<input>
<ID>IN_2</ID>96 </input>
<input>
<ID>IN_3</ID>99 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>134</ID>
<type>AI_XOR4</type>
<position>4.5,-25</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>98 </input>
<input>
<ID>IN_2</ID>96 </input>
<input>
<ID>IN_3</ID>100 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>135</ID>
<type>BE_DECODER_3x8</type>
<position>26,-14.5</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>102 </input>
<input>
<ID>IN_2</ID>101 </input>
<output>
<ID>OUT_1</ID>104 </output>
<output>
<ID>OUT_2</ID>105 </output>
<output>
<ID>OUT_3</ID>106 </output>
<output>
<ID>OUT_4</ID>107 </output>
<output>
<ID>OUT_5</ID>108 </output>
<output>
<ID>OUT_6</ID>109 </output>
<output>
<ID>OUT_7</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>136</ID>
<type>GA_LED</type>
<position>50.5,-1.5</position>
<input>
<ID>N_in0</ID>111 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>GA_LED</type>
<position>50.5,-6</position>
<input>
<ID>N_in0</ID>117 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>GA_LED</type>
<position>50.5,-10.5</position>
<input>
<ID>N_in0</ID>116 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>GA_LED</type>
<position>50.5,-15</position>
<input>
<ID>N_in0</ID>115 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>GA_LED</type>
<position>50.5,-19.5</position>
<input>
<ID>N_in0</ID>114 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>GA_LED</type>
<position>50.5,-24</position>
<input>
<ID>N_in0</ID>113 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>GA_LED</type>
<position>50.5,-28.5</position>
<input>
<ID>N_in0</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>AA_LABEL</type>
<position>-35.5,9.5</position>
<gparam>LABEL_TEXT Erorr</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-49,-2.5,-44.5,-2.5</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>-44.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-44.5,-24,-44.5,-1.5</points>
<intersection>-24 6</intersection>
<intersection>-17.5 7</intersection>
<intersection>-2.5 1</intersection>
<intersection>-1.5 8</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-44.5,-24,-43.5,-24</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>-44.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-44.5,-17.5,-43.5,-17.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>-44.5 4</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-44.5,-1.5,-21,-1.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>-44.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-49,-5,-46,-5</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>-46 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-46,-19.5,-46,-5</points>
<intersection>-19.5 11</intersection>
<intersection>-6 4</intersection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-46,-6,-21,-6</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-46 3</intersection>
<intersection>-44.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-44.5,-30.5,-44.5,-6</points>
<intersection>-30.5 6</intersection>
<intersection>-6 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-44.5,-30.5,-43.5,-30.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-44.5 5</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-46,-19.5,-43.5,-19.5</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>-46 3</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-48.5,-34.5,-48.5,-10</points>
<intersection>-34.5 6</intersection>
<intersection>-28 4</intersection>
<intersection>-21.5 9</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49,-10,-48.5,-10</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>-48.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-48.5,-28,-43.5,-28</points>
<connection>
<GID>112</GID>
<name>IN_2</name></connection>
<intersection>-48.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-48.5,-34.5,-43.5,-34.5</points>
<connection>
<GID>113</GID>
<name>IN_2</name></connection>
<intersection>-48.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-48.5,-21.5,-43.5,-21.5</points>
<connection>
<GID>111</GID>
<name>IN_2</name></connection>
<intersection>-48.5 0</intersection>
<intersection>-47 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-47,-21.5,-47,-15</points>
<intersection>-21.5 9</intersection>
<intersection>-15 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-47,-15,-21,-15</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-47 11</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-47,-32.5,-47,-7.5</points>
<intersection>-32.5 4</intersection>
<intersection>-10.5 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49,-7.5,-47,-7.5</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>-47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-47,-10.5,-21,-10.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>-47 0</intersection>
<intersection>-44 7</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-47,-32.5,-43.5,-32.5</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>-47 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-44,-26,-44,-10.5</points>
<intersection>-26 12</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>-44,-26,-43.5,-26</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>-44 7</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-3.5,-43,2</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>-3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-43,-3.5,-21,-3.5</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>-43 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-40.5,-8,-40.5,2</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-40.5,-8,-21,-8</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>-40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38,-12.5,-38,2</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-38,-12.5,-21,-12.5</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>-38 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35.5,-17,-35.5,2</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35.5,-17,-21,-17</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>-35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,-21.5,-33,2</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-33,-21.5,-21,-21.5</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>-33 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30.5,-26,-30.5,2</points>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30.5,-26,-21,-26</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>-30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-30.5,-28,2</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-28,-30.5,-21,-30.5</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>-28 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-37.5,-19.5,-21,-19.5</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<connection>
<GID>111</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36,-26,-36,-24</points>
<intersection>-26 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36,-24,-21,-24</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-37.5,-26,-36,-26</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>-36 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,-32.5,-34,-28.5</points>
<intersection>-32.5 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-28.5,-21,-28.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>-34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-37.5,-32.5,-34,-32.5</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>-34 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-15,-2.5,1.5,-2.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-15 7</intersection>
<intersection>-13.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-13.5,-12.5,-13.5,-2.5</points>
<intersection>-12.5 5</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-13.5,-12.5,1.5,-12.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>-13.5 4</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-15,-2.5,-15,-0.5</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>-2.5 1</intersection>
<intersection>-0.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-15,-0.5,39.5,-0.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>-15 7</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,-22,-11.5,-4.5</points>
<intersection>-22 4</intersection>
<intersection>-7 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11.5,-4.5,39.5,-4.5</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>-11.5 0</intersection>
<intersection>39.5 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15,-7,-11.5,-7</points>
<connection>
<GID>126</GID>
<name>OUT</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-11.5,-22,1.5,-22</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>39.5,-5,39.5,-4.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-4.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,-26,-7.5,-6.5</points>
<intersection>-26 5</intersection>
<intersection>-16 2</intersection>
<intersection>-14 3</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,-6.5,1.5,-6.5</points>
<connection>
<GID>132</GID>
<name>IN_2</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15,-16,-7.5,-16</points>
<connection>
<GID>128</GID>
<name>OUT</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-7.5,-14,39.5,-14</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>-7.5 0</intersection>
<intersection>1.5 7</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-7.5,-26,1.5,-26</points>
<connection>
<GID>134</GID>
<name>IN_2</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>1.5,-16.5,1.5,-14</points>
<connection>
<GID>133</GID>
<name>IN_2</name></connection>
<intersection>-14 3</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-20.5,-5.5,-18.5</points>
<intersection>-20.5 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5.5,-18.5,39.5,-18.5</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>-5.5 0</intersection>
<intersection>1.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-15,-20.5,-5.5,-20.5</points>
<connection>
<GID>129</GID>
<name>OUT</name></connection>
<intersection>-5.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>1.5,-18.5,1.5,-8.5</points>
<connection>
<GID>132</GID>
<name>IN_3</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-24,-9.5,-9.5</points>
<intersection>-24 4</intersection>
<intersection>-11.5 1</intersection>
<intersection>-9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,-11.5,-9.5,-11.5</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-9.5,-9.5,39.5,-9.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>-9.5 0</intersection>
<intersection>1.5 6</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-9.5,-24,1.5,-24</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>1.5,-14.5,1.5,-9.5</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>-9.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-25,-4,-23</points>
<intersection>-25 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,-25,-4,-25</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<intersection>-4 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-23,39.5,-23</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>-4 0</intersection>
<intersection>1.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>1.5,-23,1.5,-18.5</points>
<connection>
<GID>133</GID>
<name>IN_3</name></connection>
<intersection>-23 2</intersection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7,-29.5,-7,-27.5</points>
<intersection>-29.5 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-15,-29.5,-7,-29.5</points>
<connection>
<GID>131</GID>
<name>OUT</name></connection>
<intersection>-7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7,-27.5,39.5,-27.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>-7 0</intersection>
<intersection>1.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>1.5,-28,1.5,-27.5</points>
<connection>
<GID>134</GID>
<name>IN_3</name></connection>
<intersection>-27.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-16,16.5,-5.5</points>
<intersection>-16 1</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-16,23,-16</points>
<connection>
<GID>135</GID>
<name>IN_2</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-5.5,16.5,-5.5</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-17,15.5,-15.5</points>
<intersection>-17 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,-17,23,-17</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-15.5,15.5,-15.5</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-25,15.5,-18</points>
<intersection>-25 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,-18,23,-18</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-25,15.5,-25</points>
<connection>
<GID>134</GID>
<name>OUT</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-29.5,30.5,-17</points>
<intersection>-29.5 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-29.5,39.5,-29.5</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-17,30.5,-17</points>
<connection>
<GID>135</GID>
<name>OUT_1</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-25,31.5,-16</points>
<intersection>-25 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-16,31.5,-16</points>
<connection>
<GID>135</GID>
<name>OUT_2</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-25,39.5,-25</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-15,33,-11.5</points>
<intersection>-15 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-11.5,39.5,-11.5</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-15,33,-15</points>
<connection>
<GID>135</GID>
<name>OUT_3</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-20.5,34.5,-14</points>
<intersection>-20.5 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-20.5,39.5,-20.5</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-14,34.5,-14</points>
<connection>
<GID>135</GID>
<name>OUT_4</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-13,36,-7</points>
<intersection>-13 2</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-7,39.5,-7</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-13,36,-13</points>
<connection>
<GID>135</GID>
<name>OUT_5</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-12,37,-2.5</points>
<intersection>-12 2</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-2.5,39.5,-2.5</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-12,37,-12</points>
<connection>
<GID>135</GID>
<name>OUT_6</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-16,38,-11</points>
<intersection>-16 1</intersection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-16,39.5,-16</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-11,38,-11</points>
<connection>
<GID>135</GID>
<name>OUT_7</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-1.5,49.5,-1.5</points>
<connection>
<GID>136</GID>
<name>N_in0</name></connection>
<connection>
<GID>100</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-28.5,49.5,-28.5</points>
<connection>
<GID>142</GID>
<name>N_in0</name></connection>
<connection>
<GID>106</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-24,49.5,-24</points>
<connection>
<GID>141</GID>
<name>N_in0</name></connection>
<connection>
<GID>105</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-19.5,49.5,-19.5</points>
<connection>
<GID>140</GID>
<name>N_in0</name></connection>
<connection>
<GID>104</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-15,49.5,-15</points>
<connection>
<GID>139</GID>
<name>N_in0</name></connection>
<connection>
<GID>103</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-10.5,49.5,-10.5</points>
<connection>
<GID>138</GID>
<name>N_in0</name></connection>
<connection>
<GID>102</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>45.5,-6,49.5,-6</points>
<connection>
<GID>137</GID>
<name>N_in0</name></connection>
<connection>
<GID>101</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.1</PageViewport></page 9></circuit>